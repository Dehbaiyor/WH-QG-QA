�ccollections
defaultdict
q cdill._dill
_create_function
q(cdill._dill
_create_code
q(K K K KKCCt dd� �S qNh(K K K KKSCdS qNK�q))X   <ipython-input-11-f0502a42197e>qX   <lambda>qKC q))tq	Rq
X   <lambda>.<locals>.<lambda>q�qX   defaultdictq�q)hhKh))tqRqc__builtin__
__main__
hNN}qNtqRq�qRq(NN�qh h(h
c__builtin__
__main__
hNN}qNtqRq�qRq(X   WRBqG?ʻ坁>BX   WPqG?���45eX   INqG?��|���)X   JJqG?��z��cX   TOq G?i�1�P6X   NNPq!G?� 7:��,X   NNq"G?}��rlX   PRPq#G?D]��u-�X   WDTq$G?�~��c{nX   DTq%G?���=��1X   ``q&G?4�����X   PRP$q'G?$�����X   CDq(G?N���큁X   RBq)G?r��.�X   VBGq*G?vY.?�VX   NNSq+G?|B��=�_X   VBDq,G?>`:�r=X   oovq-G?J�3#�UX   JJSq.G?G ��P��X   VBZq/G?|ݠ���UX   VBPq0G?U���%Y�X   JJRq1G?$�����X   VBNq2G?A����[xX   VBq3G?a�ܟ��X   MDq4G?R���BX   CCq5G?T����X   NNPSq6G>�p�ސ�uNh�q7h h(h
c__builtin__
__main__
hNN}q8Ntq9Rq:�q;Rq<(X   VBDq=G?��n1��X   JJq>G?���J�X   RBq?G?�Z y�PX   MDq@G?��RO��X   VBZqAG?���C�ɭX   NNPqBG?k=?��%X   DTqCG?w�XK�UX   NNqDG?uk�ir�X   VBPqEG?��}}�[kX   VBqFG?��k7C�X   INqGG?s��j��X   NNSqHG?W��r�X   PRPqIG?G�XK�UX   CDqJG?0�6?s=X   VBGqKG?QU��8� X   VBNqLG?@�6?s=X   ,qMG?7�XK�UX   CCqNG?0�6?s=X   WRBqOG?#�tK��IX   oovqPG?B(�E_��X   WDTqQG?i�d�bX   TOqRG?*i�d�bX   JJRqSG?i�d�buhh=�qTh h(h
c__builtin__
__main__
hNN}qUNtqVRqW�qXRqY(X   NNPqZG?���
YX   DTq[G?�
��<�xX   PRPq\G?�i�tP��X   CDq]G?oe�d��X   NNq^G?��f�CX   VBq_G?�5fu���X   PRP$q`G?b܎��]X   NNSqaG?���5�X   JJqbG?�?�^AX   VBZqcG?>rK���X   RBqdG?�n�R\,X   JJSqeG?q�b��vX   VBGqfG?sn�R\,X   oovqgG?d��X   INqhG?Q J6��X   TOqiG?6ոH�;hX   ``qjG?h�����X   JJRqkG?NrK���X   VBNqlG?r���#�EX   NNPSqmG?g�J�&�7X   VBDqnG?>rK���X   RBSqoG?Cn�R\,X   CCqpG?.rK���X   POSqqG?6ոH�;hX   ''qrG?6ոH�;huh=hZ�qsh h(h
c__builtin__
__main__
hNN}qtNtquRqv�qwRqx(X   VBqyG?��o���X   NNqzG?�IVS/�VX   POSq{G?�1[gi�X   DTq|G?��U����X   NNPq}G?��b��:X   WRBq~G?p�KY�X   TOqG?��J���X   VBGq�G?yԓ�z4X   INq�G?�B_(�r>X   VBDq�G?��6��X   CCq�G?� )��8SX   RBq�G?�'��Ђ�X   JJq�G?�D�E�NX   RPq�G?2�@�X   .q�G?�؞�-��X   NNSq�G?����ZX   VBZq�G?D��)H�X   VBNq�G?�	�p{X�X   VBPq�G?Z�xc��?X   PRP$q�G?B�@�X   oovq�G?W7�JQX   WPq�G?2�@�X   CDq�G?lqCT�ThMG?p@���8�X   JJSq�G?D��)H�X   NNPSq�G?Y�F�kY1X   PRPq�G?g�| �X   JJRq�G?2�@�X   ``q�G?D��)H�X   RBSq�G?B�@�NG?@@���8�X   ''q�G?"�@�X   WDTq�G?"�@�X   MDq�G?Kܪ%�aMuhZhy�q�h h(h
c__builtin__
__main__
hNN}q�Ntq�Rq��q�Rq�(X   VBGq�G?�Fi���X   NNPq�G?���+��X   RPq�G?�Qs�vR%X   JJq�G?�Z�t�&X   INq�G?�=7e"Th�G?�V��ʺ�X   PRP$q�G?��8E�!�X   DTq�G?��� ��X   PRPq�G?��3�NsX   TOq�G?�Gy�%`X   NNq�G?�^��X   JJRq�G?i"$�X   VBNq�G?��>ɇjX   RBq�G?�2��y�>X   CDq�G?t���fU�X   JJSq�G?`CD���X   NNSq�G?��W
�#X   WRBq�G?rz��?�7X   VBDq�G?w��ᙆ�X   VBq�G?g��ᙆ�X   MDq�G?uo��s"X   ``q�G?l��O�X   WDTq�G?G��ᙆ�X   CCq�G?Q��i3%X   WPq�G?c8:L�mX   VBZq�G?]��Y��XX   oovq�G?a��i3%X   VBPq�G?Q��i3%X   NNPSq�G?7��ᙆ�NG?A��i3%hMG?Q��i3%X   POSq�G?7��ᙆ�uhyh��q�h h(h
c__builtin__
__main__
hNN}q�Ntq�Rq��q�Rq�(X   JJq�G?�ZZZZZZX   PRP$q�G?�X   WPq�G?�X   NNPq�G?�h�G?�������X   RBq�G?�������X   INq�G?�ddddddX   DTq�G?ť�����X   NNq�G?�xxxxxxX   TOq�G?�������X   NNSq�G?�������X   VBNq�G?�UUUUUUX   CDq�G?~X   VBq�G?�X   WRBq�G?�X   JJRq�G?�X   RPq�G?�X   VBGq�G?tX   PRPq�G?�hMG?tuh�hq�h h(h
c__builtin__
__main__
hNN}q�Ntq�Rqׅq�Rq�(h�G?�����X   NNq�G?�.����X   NNSq�G?�S#eX   INq�G?�WAh�JX   TOq�G?�f���\X   JJq�G?�S#eX   CCq�G?����X   NNPq�G?������X   VBNq�G?��pŎg�X   VBZq�G?s�pŎg�hMG?s�pŎg�X   RBq�G?zWAh�JX   WPq�G?zWAh�JX   JJSq�G?jWAh�JX   NNPSq�G?jWAh�JX   JJRq�G?s�pŎg�X   VBDq�G?jWAh�JX   VBGq�G?s�pŎg�X   ''q�G?jWAh�JX   VBq�G?jWAh�Juh�h��q�h h(h
c__builtin__
__main__
hNN}q�Ntq�Rq�q�Rq�(NG?�)����X   ``q�G?bN_��X   VBDq�G?RN_��h�G?[u�M�܈X   ''q�G?y+�\c�'X   WPq�G?RN_��X   oovq�G?RN_��uh�N�q�h h(h
c__builtin__
__main__
hNN}q�Ntq�Rq��q�Rq�NG?�      sNh�q�h h(h
c__builtin__
__main__
hNN}q�Ntq�Rr   �r  Rr  (X   NNSr  G?�[�6���X   NNr  G?���e8�RX   VBDr  G?�.��_X   VBZr  G?ќ@�P�X   JJRr  G?*,�����X   JJr  G?���?%X   NNPr	  G?�7+�p�|X   RBr
  G?>�S�`X   MDr  G?�Q��T_KX   VBPr  G?��/����X   INr  G?UDQࡠ�X   VBGr  G?\w@ZMkX   CDr  G?���AZ�X   VBr  G?Oh�s%��hMG?At����X   PRPr  G?$���;�X   oovr  G?,�����X   JJSr  G?,�����X   WRBr  G?h�s%��X   ``r  G?,��~�[X   TOr  G?���;�X   WPr  G?���;�X   VBNr  G?'���\cbX   DTr  G?>�yFX   WDTr  G?���;�X   NNPSr  G?h�s%��X   RBSr  G?���;�uhj  �r  h h(h
c__builtin__
__main__
hNN}r  Ntr  Rr   �r!  Rr"  (X   VBDr#  G?�B^З�&X   INr$  G?�8�8�X   VBPr%  G?�O)�X   MDr&  G?�O)�h�G?���<X   VBZr'  G?�O)�X   NNr(  G?��%�	{BX   WPr)  G?YH�����X   CCr*  G?iH�����X   JJr+  G?o��<�XX   DTr,  G?��<�X~X   NNSr-  G?�a�����X   WRBr.  G?b����/hX   RBr/  G?iH�����X   TOr0  G?iH�����hMG?iH�����X   VBGr1  G?YH�����X   VBr2  G?YH�����X   VBNr3  G?|q�q�NG?YH�����X   RPr4  G?YH�����X   POSr5  G?o��<�XX   NNPr6  G?iH�����uj  j#  �r7  h h(h
c__builtin__
__main__
hNN}r8  Ntr9  Rr:  �r;  Rr<  (X   NNPr=  G?�G���pX   PRP$r>  G?z(젹HX   INr?  G?��V[u�6X   PRPr@  G?���R>�fX   ``rA  G?Y]���k�X   DTrB  G?�~W�ůX   VBNrC  G?șdT:%X   WDTrD  G?d�]W���X   JJrE  G?���Ho`�X   NNSrF  G?��0�C�pX   TOrG  G?������X   NNrH  G?��-	]1�h�G?��t����X   VBGrI  G?�nI�ȂgX   RBrJ  G?�r��.��X   WPrK  G?�b��H�{X   oovrL  G?t�]W���X   CDrM  G?l��R>�fX   RPrN  G?���ڤ��X   VBDrO  G?d�]W���X   VBrP  G?j�܆���X   JJSrQ  G?Y]���k�X   WRBrR  G?d�]W���X   JJRrS  G?f2=#�lX   RBSrT  G?Y]���k�hMG?V2=#�lX   CCrU  G?c}�)��X   NNPSrV  G?S}�)��NG?V2=#�lX   VBZrW  G?9]���k�X   ''rX  G?9]���k�uj=  hz�rY  h h(h
c__builtin__
__main__
hNN}rZ  Ntr[  Rr\  �r]  Rr^  (X   INr_  G?��mb̐X   VBDr`  G?��tY�Xh�G?�|���<X   TOra  G?�SV1>)�X   NNPrb  G?��� %X   DTrc  G?�P!�H�LX   ''rd  G?U,x��hMG?�/��X   MDre  G?vpE��X   NNrf  G?���cdXX   NNSrg  G?�ԉĺ>�X   PRP$rh  G?bc@v ��X   CCri  G?�/��X   RPrj  G?O4LV:(X   POSrk  G?y��оX   VBZrl  G?������X   WDTrm  G?}�!��-�X   VBrn  G?{��0�DX   RBro  G?������X   VBGrp  G?x˨a;`�X   VBPrq  G?�&Hx�mX   VBNrr  G?�ώ�D�X   JJrs  G?z0D�6bX   WRBrt  G?gg9@��X   WPru  G?\�|�+&X   PRPrv  G?lj��`�eX   oovrw  G?Z��f �#X   CDrx  G?bc@v ��NG?e,x��X   ``ry  G?[�3�!�X   JJRrz  G?Aԛ�U�X   NNPSr{  G?6I��NX   JJSr|  G?1ԛ�U�X   RBSr}  G?6I��Nuhzj_  �r~  h h(h
c__builtin__
__main__
hNN}r  Ntr�  Rr�  �r�  Rr�  (X   WRBr�  G?g�љX   PRP$r�  G?�pd���X   NNPr�  G?��<�X~X   NNr�  G?������OX   CDr�  G?�FR�8th�G?������X   WPr�  G?�c{��9�X   WDTr�  G?�\"q
kjX   PRPr�  G?w� 0�4�X   DTr�  G?Ӕy�o��X   INr�  G?����X�X   JJSr�  G?Z�b�D�X   VBGr�  G?�:�i��MX   NNSr�  G?���_���X   JJr�  G?���tX   RBr�  G?cՄ��f�X   oovr�  G?R���rX   TOr�  G?U̱���X   ``r�  G?oEf�S�X   VBNr�  G?`B�I��hMG?A�W0�;X   JJRr�  G?W�!ϸ�X   VBDr�  G?@pd���X   NNPSr�  G?T^�pVNX   CCr�  G?DB�,^�X   MDr�  G?!']���lX   VBZr�  G?F�'�{��X   VBPr�  G?']���lX   VBr�  G?']���lX   RBSr�  G?�'�{��NG?5q5M�Guj_  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   PRPr�  G?�g�$��X   JJr�  G?�p�S�h�G?�D�#pbX   NNr�  G?~���E�X   TOr�  G?�VL���X   VBGr�  G?��ڥ��X   NNPr�  G?����{AX   INr�  G?��ڥ��X   VBZr�  G?��ڥ��X   VBDr�  G?�Ik:�1X   RBr�  G?���<�BX   NNSr�  G?��ڥ��X   VBNr�  G?����E�X   DTr�  G?���N�X   MDr�  G?y��N�X   VBPr�  G?��O��AX   CCr�  G?d�ڥ��X   VBr�  G?y��N�hMG?d�ڥ��X   oovr�  G?d�ڥ��X   PRP$r�  G?d�ڥ��X   WPr�  G?d�ڥ��uj�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   VBDr�  G?�M�"6�X   VBZr�  G?���-�ɟX   VBPr�  G?�b^8X   RBr�  G?���K�X   MDr�  G?�S�=�X   VBr�  G?s�"�f�X   WDTr�  G?s�"�f�h�G?}S�=�uj�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   VBGr�  G?�4YZ;<X   DTr�  G?�0q�;�X   PRPr�  G?���_��X   NNPr�  G?�AoZ��X   RBr�  G?�
��3�X   INr�  G?��)�[&XX   VBNr�  G?áh�6�X   TOr�  G?������X   JJr�  G?��cjM�h�G?�EV���X   ''r�  G?f
��3�X   NNSr�  G?�
��3�X   PRP$r�  G?�tg�bX   CDr�  G?���_��X   RPr�  G?�9��t- X   NNr�  G?�^"p���X   WRBr�  G?��Q�F|X   ``r�  G?r^"p���X   VBr�  G?mcjM���X   oovr�  G?���˦�hMG?y���4X   WPr�  G?r^"p���X   VBDr�  G?f
��3�X   WDTr�  G?]cjM���X   CCr�  G?mcjM���X   JJRr�  G?f
��3�X   VBPr�  G?]cjM���X   MDr�  G?]cjM���uj�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   RPr�  G?��?��X   NNPr�  G?�.��f�X   DTr�  G?���5�KX   RBr�  G?�>���X   NNSr�  G?�ɕ�{��X   INr�  G?�.��f�h�G?�b�O��X   NNr�  G?�5-�*^X   JJr�  G?����V(fhMG?�ɕ�{��X   VBNr�  G?��P�x_�X   VBr�  G?�}R	��X   ``r�  G?zb�O��X   TOr�  G?�#s�Ʋ�X   PRPr�  G?��?��X   POSr�  G?�b�O��X   JJRr�  G?�}R	��X   oovr�  G?�}R	��X   VBDr�  G?sɕ�{��X   PRP$r�  G?��?��X   WRBr�  G?�}R	��X   WPr   G?�}R	��X   CCr  G?�ɕ�{��X   VBGr  G?�b�O��X   JJSr  G?jb�O��X   VBZr  G?jb�O��X   VBPr  G?jb�O��X   ''r  G?jb�O��X   CDr  G?jb�O��X   WDTr  G?jb�O��uj�  j�  �r	  h h(h
c__builtin__
__main__
hNN}r
  Ntr  Rr  �r  Rr  (h�G?�X   INr  G?�������X   NNr  G?�X   TOr  G?�������X   WPr  G?�X   NNSr  G?�������X   JJr  G?�X   RBr  G?�X   NNPr  G?�X   DTr  G?�X   ''r  G?�X   PRP$r  G?�X   oovr  G?�hMG?�X   CCr  G?�X   VBNr  G?�X   WRBr  G?�uj�  h��r  h h(h
c__builtin__
__main__
hNN}r  Ntr   Rr!  �r"  Rr#  NG?�      sX   VBr$  h��r%  h h(h
c__builtin__
__main__
hNN}r&  Ntr'  Rr(  �r)  Rr*  (X   POSr+  G?��[}���X   NNr,  G?�yf톙X   NNPr-  G?�H#0b�zh�G?��IfQX   INr.  G?����NG?\&�9.�X   NNSr/  G?�Z��PX   VBGr0  G?x�ޒ�X   CCr1  G?�� ���X   VBr2  G?��s>u�X   TOr3  G?��s>u�X   RBr4  G?�dI囶hMG?|&�9.�X   DTr5  G?��s>u�X   ''r6  G?l&�9.�X   ``r7  G?\&�9.�X   MDr8  G?q�1C�$X   VBDr9  G?�Z��PX   NNPSr:  G?q�1C�$X   JJr;  G?����X   CDr<  G?����X   oovr=  G?q�1C�$X   VBNr>  G?�Z��PX   VBZr?  G?e���X   PRP$r@  G?q�1C�$X   JJSrA  G?\&�9.�X   PRPrB  G?\&�9.�X   VBPrC  G?\&�9.�X   WPrD  G?\&�9.�uh�j+  �rE  h h(h
c__builtin__
__main__
hNN}rF  NtrG  RrH  �rI  RrJ  (X   NNPrK  G?���B�X   NNrL  G?���ټ�MX   JJrM  G?���ѹ{X   JJRrN  G?b�U1�x�X   VBGrO  G?q �ڼ�X   NNPSrP  G?1�nM&GX   NNSrQ  G?��+�%��X   ``rR  G?yj����vX   RBSrS  G?q �ڼ�X   JJSrT  G?�-����X   CDrU  G?�����X   CCrV  G?`��hS��X   VBNrW  G?���cH�^h�G?���E{uX   VBDrX  G?k��X��^X   WPrY  G?:��s�"�X   INrZ  G?q �ڼ�X   DTr[  G?q �ڼ�X   PRPr\  G?A�nM&GX   VBPr]  G?\�s=]��hMG?J��s�"�X   VBZr^  G?Z��s�"�X   RBr_  G?c�<��/X   RPr`  G?1�nM&GX   VBra  G?F	�o�X   MDrb  G?:��s�"�X   WDTrc  G?1�nM&GX   PRP$rd  G?1�nM&GX   TOre  G?1�nM&Guj+  jK  �rf  h h(h
c__builtin__
__main__
hNN}rg  Ntrh  Rri  �rj  Rrk  (X   CCrl  G?�l�M��X   NNrm  G?Ņ��XZ�h�G?�/�A��X   VBPrn  G?��Q���hMG?�A��40X   INro  G?��c�qFX   POSrp  G?�ɠ�|�X   VBrq  G?��Q���X   VBDrr  G?���=+TX   MDrs  G?k/�A��4X   NNPrt  G?�1�8�tX   NNSru  G?��ɠ�}X   CDrv  G?���	��X   DTrw  G?b��!�xX   VBZrx  G?�Q����X   RBry  G?��Q���X   ''rz  G?��Q���X   NNPSr{  G?�/�A��4X   VBGr|  G?k/�A��4X   TOr}  G?r��!�xX   VBNr~  G?���!�xX   WDTr  G?b��!�xX   JJr�  G?v��ajzVX   WPr�  G?b��!�xNG?b��!�xX   oovr�  G?b��!�xX   PRP$r�  G?b��!�xX   ``r�  G?r��!�xujK  jl  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   VBr�  G?���M�,�X   NNPr�  G?��^NhlfX   PRP$r�  G?���@X   NNr�  G?���ہ� X   DTr�  G?��Z�)_6X   INr�  G?j��@X   WDTr�  G?����X   NNSr�  G?������X   WPr�  G?�J��A��X   CDr�  G?z��@X   VBZr�  G?w�8r X   JJr�  G?�T�*�5LX   PRPr�  G?aW���X   VBDr�  G?���@X   VBNr�  G?l���΀X   RBr�  G?���A80X   NNPSr�  G?z��@X   VBGr�  G?W�8r X   VBPr�  G?W�8r X   WRBr�  G?g�8r h�G?G�8r X   oovr�  G?aW���X   JJSr�  G?G�8r X   TOr�  G?G�8r ujl  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   DTr�  G?�\(��X   NNr�  G?�z�G�{X   PRP$r�  G?��Q��X   WPr�  G?�p��
=qh�G?���
=p�X   NNSr�  G?�\(��X   NNPr�  G?��Q��X   INr�  G?�
=p��
X   JJRr�  G?�z�G�{X   JJr�  G?�\(��X   RPr�  G?�z�G�{X   PRPr�  G?�
=p��
X   RBr�  G?���
=p�X   CCr�  G?�z�G�{X   VBDr�  G?tz�G�{X   ''r�  G?tz�G�{X   TOr�  G?�z�G�{X   VBNr�  G?�������X   CDr�  G?�z�G�{X   VBGr�  G?~�Q��X   JJSr�  G?tz�G�{X   VBZr�  G?tz�G�{hMG?�z�G�{X   oovr�  G?tz�G�{X   WRBr�  G?tz�G�{X   VBr�  G?tz�G�{X   ``r�  G?~�Q��uj�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   JJr�  G?�x���X   NNr�  G?�e�>{:$X   NNSr�  G?�A���RX   NNPr�  G?�_u'X   PRPr�  G?DӾ&.�X   JJSr�  G?�9FJ�iX   RBSr�  G?z��/��X   VBDr�  G?s�� ���X   JJRr�  G?z��/��X   NNPSr�  G?s�� ���X   VBGr�  G?xL]��6�X   CDr�  G?���z[��X   VBZr�  G?m�M;��cX   INr�  G?}�M;��cX   VBNr�  G?cn5ͪ�X   VBr�  G?cn5ͪ�X   VBPr�  G?DӾ&.�X   WPr�  G?[��e�>{X   RBr�  G?j��/��X   ``r�  G?s�� ���X   DTr�  G?a[_u'X   oovr�  G?j��/��X   TOr�  G?;��e�>{h�G?a[_u'hMG?DӾ&.�X   WRBr�  G?;��e�>{X   MDr�  G?TӾ&.�X   PRP$r�  G?K��e�>{X   CCr�  G?;��e�>{uj�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   NNr�  G?�Q��BX   JJr�  G?�g��t�hMG?g׈��X   VBNr�  G?x��� �*X   INr�  G?�XmF��4X   NNPr�  G?�sI9��X   NNSr�  G?��,4��X   CDr�  G?�n��|iX   VBGr�  G?i��wM�h�G?�d '��nX   ``r�  G?_�
���X   MDr�  G?*���ҞX   TOr�  G?x�:�+��X   CCr�  G?���+��X   VBDr�  G?]G��N]X   JJSr�  G?p�.y�X   WPr�  G?Rg{���X   RBSr�  G?XB�i
V�X   RBr�  G?`P�c�XX   VBZr�  G?Wls���JX   RPr�  G?$��+��X   ''r�  G?7ls���JX   DTr�  G?@�.y�X   WRBr�  G?4��+��X   WDTr�  G?E�"L�� X   VBPr�  G?\qg����X   oovr   G?D��+��X   POSr  G?Bg{���X   NNPSr  G?^�VA��X   VBr  G?J���ҞX   PRPr  G?$��+��X   JJRr  G?4��+��NG?$��+��uj�  j�  �r  h h(h
c__builtin__
__main__
hNN}r  Ntr  Rr	  �r
  Rr  (h�G?��b1��GX   NNPr  G?�y!�BBX   NNr  G?�%�R	�YX   VBDr  G?�X��@�X   INr  G?�g�x��X   TOr  G?����H[�X   VBNr  G?���A�,ihMG?�$����X   ``r  G?[DD�-הX   VBGr  G?}O�G�X   CDr  G?T���X   WDTr  G?���+��7X   WRBr  G?b�b����X   NNSr  G?�kThX   POSr  G?t�ai�X   PRP$r  G?5�7$�vX   VBZr  G?�%��x
�X   RBr  G?���%�9X   CCr  G?�-����X   ''r  G?t���vD�X   VBr  G?y[�m�}X   JJr  G?8hnn�X   PRPr   G?R��7���X   DTr!  G?r�Isu�X   VBPr"  G?����vD�X   MDr#  G?�\)O�YX   WPr$  G?eD�
(&X   RPr%  G?*-����X   JJRr&  G?5�7$�vX   oovr'  G?T-f%��NG?P��I6�X   JJSr(  G?.����rX   RBSr)  G?1s_CP��X   NNPSr*  G?s_CP��uj�  h��r+  h h(h
c__builtin__
__main__
hNN}r,  Ntr-  Rr.  �r/  Rr0  (NG?��]t��X   ''r1  G?]�3���X   ``r2  G?B�Rj�%uh�G?B�Rj�%uX   VBr3  G? �IBB��X   CCr4  G?�m�d1�X   WPr5  G? �IBB��X   WDTr6  G?�IBB��X   WRBr7  G?�m�d1�X   oovr8  G?$�[��~�X   NNr9  G? �IBB��X   VBDr:  G? �IBB��X   JJr;  G?�IBB��X   RBr<  G?�IBB��X   INr=  G?(�m�d1�X   NNPr>  G? �IBB��X   PRPr?  G? �IBB��X   DTr@  G?�m�d1�uNh�rA  h h(h
c__builtin__
__main__
hNN}rB  NtrC  RrD  �rE  RrF  (X   WPrG  G?���ZhX   WDTrH  G?��t���X   PRP$rI  G?vx�OX   VBGrJ  G?����^�X   CDrK  G?��ecW�MX   JJrL  G?���Ӵ�X   oovrM  G?xT�A�$qX   NNPrN  G?�� O��X   INrO  G?�=(�]&X   NNrP  G?��QW��yX   DTrQ  G?��>�yvX   WRBrR  G?�Xr�6�X   RBrS  G?g �����X   PRPrT  G?vx�OX   VBNrU  G?`�y�p+�X   NNSrV  G?�z��`�X   JJSrW  G?X���3X   JJRrX  G?U;�^r�X   VBDrY  G?A���
IX   ``rZ  G?A���
IX   NNPSr[  G?,O��C�hMG?,O��C�X   RPr\  G?,O��C�X   VBr]  G?,O��C�X   CCr^  G?,O��C�uhjG  �r_  h h(h
c__builtin__
__main__
hNN}r`  Ntra  Rrb  �rc  Rrd  (X   NNre  G?�j�%X   NNPrf  G?��y=�q[X   JJrg  G?�o��k�h�G?�|6du)X   INrh  G?����8��X   POSri  G?G��� X   VBZrj  G?���fXX   TOrk  G?W��� X   NNSrl  G?��`XX   VBDrm  G?�o(��'X   VBPrn  G?p�N��"X   MDro  G?b��P��X   VBGrp  G?fÈ���X   DTrq  G?S�k�dUX   JJRrr  G?U�)�k;+X   PRPrs  G?S�k�dUX   CDrt  G?����T@X   WPru  G??��vmmVX   ''rv  G??��vmmVX   RBrw  G?aЭ����X   WRBrx  G?QЭ����hMG?S�k�dUX   WDTry  G?7��� X   CCrz  G?/��vmmVX   ``r{  G?7��� X   oovr|  G?7��� NG?/��vmmVX   VBr}  G?7��� X   JJSr~  G?7��� ujG  je  �r  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   CCr�  G?p2��6X   VBDr�  G?�����-X   VBGr�  G?[�zc�+�X   VBNr�  G?n�j2��h�G?�0H���X   INr�  G?�Y����'X   NNr�  G?��a�&K'X   POSr�  G?~n>�:hMG?`��H9�X   VBZr�  G?��b��FX   NNSr�  G?�o!ݳ� X   VBPr�  G?��\L��IX   TOr�  G?d���G�X   RBr�  G?{_�gD�X   NNPr�  G?P��H9�X   MDr�  G?�P��
T�X   DTr�  G?I��lV[X   RBSr�  G?$��V�|X   JJr�  G?`L��kUX   CDr�  G?:�~ps�PX   WRBr�  G?>n>�:X   WDTr�  G?LkvWz�EX   PRPr�  G?*�~ps�PX   VBr�  G?$��V�|X   ''r�  G?$��V�|X   oovr�  G?$��V�|X   WPr�  G?0��H9�NG?$��V�|X   JJRr�  G?*�~ps�PX   JJSr�  G?�~ps�PX   ``r�  G?�~ps�Puje  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   NNr�  G?ߌ��-�X   VBr�  G?��ғ_D�X   RBr�  G?�gb���X   VBDr�  G?�2ĳ�TEX   NNPr�  G?�x����X   DTr�  G?�/���X   JJr�  G?�͊9���X   NNSr�  G?��G87�X   VBNr�  G?�quB��=X   PRP$r�  G?}�D�X   JJRr�  G?��ғ_D�X   VBZr�  G?�`K���iX   WPr�  G?��*��iX   CDr�  G?}�D�X   WDTr�  G?m�D�X   INr�  G?��/���X   VBGr�  G?��Y�<��X   TOr�  G?ZO"P��X   PRPr�  G?`quB��=X   JJSr�  G?g=���"X   WRBr�  G?pquB��=X   VBPr�  G?pquB��=X   MDr�  G?g=���"NG?JO"P��X   CCr�  G?c�Y�<��X   ``r�  G?JO"P��X   POSr�  G?JO"P��h�G?S�Y�<��X   RBSr�  G?S�Y�<��hMG?JO"P��uj�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   VBDr�  G?���S�QX   INr�  G?�S���q9h�G?��ƴ�.X   NNr�  G?��R����X   MDr�  G?�	����X   VBPr�  G?�n�5Ζ�X   NNSr�  G?�ļ�C%"X   VBNr�  G?��.���X   CDr�  G?Sf����X   VBZr�  G?���x�hMG?��P�{`�X   CCr�  G?�@C�$�3X   DTr�  G?x@C�$�3X   TOr�  G?�ў�U�X   WPr�  G?cf����X   ''r�  G?sf����X   RBr�  G?�@C�$�3X   WRBr�  G?]�_�X   NNPr�  G?z�~A��X   JJr�  G?�f����X   WDTr�  G?x@C�$�3X   VBGr�  G?m�_�X   POSr�  G?p��!��
X   VBr�  G?p��!��
X   PRP$r�  G?Sf����X   oovr�  G?��I�hHX   RBSr�  G?Sf����uj�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   NNPr�  G?�g3�&$X   PRPr�  G?�+c�4X   PRP$r�  G?zm��mX   NNr�  G?��ڭ7�,X   DTr�  G?�N6]CX   INr�  G?�����X   VBNr�  G?�S0ڑ�X   oovr�  G?u=K~�wUX   WDTr�  G?\��Y;�X   WRBr�  G?a�'dI
�X   RPr�  G?u|����X   NNSr�  G?����87X   TOr�  G?�7b�)X   WPr�  G?sF�\Vh�G?�we��X   CDr�  G?w���$X   JJr�  G?�DQp;�X   VBGr�  G?�I���X   RBr�  G?�P�D��X   ``r�  G?e��^ bKX   JJRr�  G?e��^ bKX   VBr�  G?l'��P�X   JJSr�  G?b�"���X   CCr�  G?V���87X   RBSr�  G?T�؟��_X   VBZr�  G?;� ��e�hMG?I�UW���X   VBDr   G?O��κ��X   NNPSr  G?R�"���X   VBPr  G?��κ��NG?E��^ bKX   MDr  G?'���$X   ''r  G?��κ��X   POSr  G?��κ��uX   VBr  h��r  h h(h
c__builtin__
__main__
hNN}r  Ntr	  Rr
  �r  Rr  (h�G?ȹEz�*X   INr  G?����XX   VBGr  G?�FI۲cX   DTr  G?���efX   NNr  G?�D9��X   TOr  G?��s+02X   NNSr  G?��s+02X   NNPr  G?�K�f�~oX   PRP$r  G?�I۲b�X   WPr  G?�	c�Q��X   CCr  G?�	c�Q��X   WRBr  G?�D9��X   JJr  G?�	c�Q��X   ''r  G?t��efX   CDr  G?~D9��X   RBr  G?���v옹X   JJSr  G?~D9��X   WDTr  G?~D9��X   JJRr  G?~D9��X   PRPr  G?t��efX   oovr   G?t��efhMG?t��efX   VBNr!  G?t��efX   ``r"  G?~D9��uX   INr#  jH  �r$  h h(h
c__builtin__
__main__
hNN}r%  Ntr&  Rr'  �r(  Rr)  (X   NNr*  G?��Ռ8�_X   NNSr+  G?�9��f�X   JJr,  G?��;-n�X   CDr-  G?�K�Ew�`X   NNPr.  G?�K�Ew�`X   VBDr/  G?��?	ITX   PRPr0  G?�ލ���mX   DTr1  G?��7Q��X   VBZr2  G?|M/�ގX   INr3  G?�'� )*tX   oovr4  G?d�9��gX   VBPr5  G?|M/�ގX   VBGr6  G?n��Ռ8�X   RBr7  G?n��Ռ8�X   WPr8  G?d�9��gX   JJRr9  G?^��Ռ8�X   NNPSr:  G?T�9��gX   JJSr;  G?T�9��gX   RPr<  G?T�9��gX   TOr=  G?T�9��gujH  j*  �r>  h h(h
c__builtin__
__main__
hNN}r?  Ntr@  RrA  �rB  RrC  (X   VBDrD  G?��M�X   INrE  G?c��~�hMG?:9栰�X   POSrF  G?�k�l���h�G?��eЂGX   NNrG  G?���`�iX   RBrH  G?�7Lq3�X   CCrI  G?z���>!X   WDTrJ  G?o:9栰�X   VBZrK  G?�_Ob��X   TOrL  G?��{��NX   VBPrM  G?�F�H6��X   JJrN  G?_:9栰�X   NNSrO  G?�R�̚�X   VBGrP  G?r7Lq3�X   CDrQ  G?d�{��NX   NNPrR  G?r7Lq3�X   VBNrS  G?t�{��NX   MDrT  G?�*���X   DTrU  G?d�{��NX   WPrV  G?T�{��NX   JJRrW  G?T�{��NX   oovrX  G?T�{��NX   WRBrY  G?T�{��NuX   VBrZ  h��r[  h h(h
c__builtin__
__main__
hNN}r\  Ntr]  Rr^  �r_  Rr`  (h�G?��CB�-hX   TOra  G?�e����X   NNSrb  G?���M�X   NNrc  G?�=)�I��X   INrd  G?�,��y��X   NNPre  G?�C�
U��X   oovrf  G?`C�
U��X   ''rg  G?k���6�X   WPrh  G?pC�
U��X   JJri  G?���c��X   CCrj  G?�%��X   NNPSrk  G?e��c��X   VBrl  G?�����gYX   VBNrm  G?pC�
U��X   RBrn  G?���6�Y�X   CDro  G?e��c��hMG?xe�����X   DTrp  G?u��c��X   VBGrq  G?u��c��X   WRBrr  G?k���6�X   PRPrs  G?e��c��NG?U��c��X   JJRrt  G?U��c��X   POSru  G?U��c��X   VBZrv  G?U��c��X   ``rw  G?U��c��uX   WPrx  jf  �ry  h h(h
c__builtin__
__main__
hNN}rz  Ntr{  Rr|  �r}  Rr~  (X   CCr  G?mn��4m%X   NNr�  G?�n��4m%X   NNPr�  G?��ɻ��X   VBDr�  G?��* ���X   NNSr�  G?�L�	�X   NNPSr�  G?��ɻ��X   POSr�  G?�+:�ޕ X   VBZr�  G?�%gQ��h�G?�n��4m%X   INr�  G?�+:�ޕ X   JJr�  G?�%gQ�X   RBr�  G?}n��4m%X   VBNr�  G?mn��4m%X   VBPr�  G?��ɻ��X   VBGr�  G?x���JX   MDr�  G?mn��4m%hMG?c�Z"�nX   CDr�  G?mn��4m%uj  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   NNr�  G?����ÙX   NNPr�  G?ѥޘQ�AX   INr�  G?����j3�X   VBGr�  G?r}�a��X   VBDr�  G?�~j�X   CDr�  G?z�_bO�X   VBr�  G?�ٍ��hMG?�x��zFbh�G?���}m$�X   ''r�  G?y6k�*�X   TOr�  G?�1Db��X   RBr�  G?�c*�h�X   NNSr�  G?�-a`�c�X   VBPr�  G?�N��ЅX   JJr�  G?y6k�*�X   POSr�  G?�A�9�nX   MDr�  G?pλ�Aq�X   WRBr�  G?J�_bO�X   VBNr�  G?��ޘQ�AX   DTr�  G?~@�NB��X   CCr�  G?�λ�Aq�X   VBZr�  G?��ޘQ�AX   oovr�  G?w��u��NG?Z�_bO�X   NNPSr�  G?y6k�*�X   WPr�  G?T+G����X   WDTr�  G?T+G����uj`  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   DTr�  G?��N���KX   JJr�  G?�H�v>�tX   NNr�  G?���^/X   VBr�  G?��'���.X   INr�  G?�S�,���X   VBDr�  G?è�R�xX   CCr�  G?l`���9�X   NNPr�  G?�H�v>�tX   VBZr�  G?���_�X   RBr�  G?������6X   TOr�  G?�ɛ}�CfX   RPr�  G?|`���9�X   VBGr�  G?�H�v>�tX   VBPr�  G?�2A�L�h�G?�p�}V��X   VBNr�  G?��_�>X   ``r�  G?�H�v>�tX   MDr�  G?���4�r�X   WDTr�  G?b�N���KX   oovr�  G?l`���9�X   PRP$r�  G?b�N���KX   WRBr�  G?r�N���KhMG?l`���9�X   NNSr�  G?r�N���KX   WPr�  G?l`���9�X   JJSr�  G?b�N���KX   JJRr�  G?l`���9�X   POSr�  G?b�N���KX   CDr�  G?b�N���Kuj�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   NNr�  G?���/X   ''r�  G?���/9h�G?���/9X   JJr�  G?��Ƈ�4?X   JJSr�  G?�X��Ƈ�X   JJRr�  G?���/9X   WPr�  G?���/9X   NNSr�  G?�X��Ƈ�X   VBPr�  G?���/9X   RBr�  G?���/9X   NNPr�  G?������X   INr�  G?���/9X   VBDr�  G?���/9X   RBSr�  G?�X��ƈX   ``r�  G?���/9hMG?���/9uj�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   NNr�  G?�wg&�auX   VBNr�  G?�sΡ�TX   INr�  G?�"����h�G?�:��,�`X   CCr�  G?���
��dX   ``r�  G?�wp��X   NNPr�  G?�R�D�hMG?���DuNX   NNSr�  G?��b(	�dX   TOr�  G?��M��X   VBDr�  G?��؞�uX   POSr�  G?�g�}H!8X   JJr�  G?��shYX   PRPr�  G?c�ȼw �X   VBr�  G?~���D��X   VBGr�  G?�a|Z���X   DTr�  G?wf��"F-X   VBZr�  G?��# x�X   VBPr�  G?���.�NX   WDTr�  G?��|��X   oovr�  G?RC��R�X   WPr�  G?p��!�S"X   WRBr�  G?pR��˻�X   RBr�  G?�J�m|iNX   ''r�  G?Ke~��k"X   RBSr�  G?=9˷�X   MDr   G?w�#Ź� X   CDr  G?fԔW'��X   JJRr  G?-9˷�X   RPr  G?@p�s{X   PRP$r  G?9˷�X   NNPSr  G?0p�s{NG?UZl0 X   JJSr  G?"C��R�uj�  j�  �r  h h(h
c__builtin__
__main__
hNN}r  Ntr	  Rr
  �r  Rr  (h�G?� ���IhMG?�(���xX   VBDr  G?�)F����X   VBNr  G?�%TC�{yX   INr  G?��^�&L�X   NNr  G?��H@�f�X   TOr  G?��wxDvX   RBr  G?�����X   CCr  G?��4l�X�X   VBPr  G?�����\lX   NNSr  G?���U�UX   WDTr  G?���4�KNX   VBr  G?��"BÊ�X   oovr  G?Z����\lX   VBZr  G?��>N�cX   ''r  G?pƘnf:1X   JJr  G?��Q�X   NNPr  G?�ΉBQ�X   VBGr  G?z&�3�Z�X   PRPr  G?]����f�X   CDr  G?Z����\lX   JJRr   G?G��P�R'X   WPr!  G?R�׊rA	X   DTr"  G?�Ƙnf:1X   MDr#  G?}����f�X   POSr$  G?h��ޖU�NG?l�O�a�X   WRBr%  G?o����m�X   PRP$r&  G?I�4l�X�X   RPr'  G?A�7�l=�X   RBSr(  G?E��4�KNX   ``r)  G?\��cDX   JJSr*  G?/����m�X   NNPSr+  G?����m�uj�  j�  �r,  h h(h
c__builtin__
__main__
hNN}r-  Ntr.  Rr/  �r0  Rr1  (X   DTr2  G?�0ѐX   CDr3  G?�0ѐX   NNr4  G?�Cީ=�X   JJr5  G?�\�����X   NNSr6  G?�Cީ=�h�G?�0ѐX   INr7  G?s0ѐX   NNPr8  G?��u�
�^X   VBNr9  G?s0ѐX   ``r:  G?s0ѐX   TOr;  G?s0ѐX   ''r<  G?s0ѐX   JJSr=  G?��_A}�uj�  j2  �r>  h h(h
c__builtin__
__main__
hNN}r?  Ntr@  RrA  �rB  RrC  (X   NNrD  G?�UUUUUUX   RBSrE  G?�UUUUUUX   JJrF  G?ڪ�����X   NNPrG  G?�      ujD  j�  �rH  h h(h
c__builtin__
__main__
hNN}rI  NtrJ  RrK  �rL  RrM  (X   NNrN  G?���Zj��X   NNPrO  G?�& �LA]X   INrP  G?ܜ�:�Vh�G?�A\���1X   WPrQ  G?t����� X   TOrR  G?�_�#��{X   WRBrS  G?s��Zj��X   PRPrT  G?J%	��5X   RBrU  G?���1rbX   DTrV  G?�>�H��X   RPrW  G?�W& �LAX   VBNrX  G?�;�6w�mX   VBDrY  G?Qn�BsyX   ``rZ  G?qn�BsyX   WDTr[  G?g�H��^�X   JJr\  G?��;�6xX   oovr]  G?Qn�BsyX   NNSr^  G?{;�6w�mX   NNPSr_  G?An�BsyX   VBZr`  G?J%	��5X   VBGra  G?eɈ+�WhMG?eɈ+�WX   JJSrb  G?Qn�BsyX   CCrc  G?g�H��^�X   VBPrd  G?An�BsyX   JJRre  G?An�BsyX   CDrf  G?UɈ+�WX   ''rg  G?An�BsyX   PRP$rh  G?An�BsyX   MDri  G?An�Bsyuj�  jN  �rj  h h(h
c__builtin__
__main__
hNN}rk  Ntrl  Rrm  �rn  Rro  (h�G?�՟��5X   INrp  G?���B-GX   CCrq  G?�8N��X   NNrr  G?��B-Gf�X   VBGrs  G?�8N��X   VBDrt  G?�j;5��[X   NNSru  G?�b�O�BX   VBNrv  G?�b�O�BX   WDTrw  G?�8N��X   RBrx  G?w8N��X   TOry  G?�����D�X   CDrz  G?b�r[��X   DTr{  G?��r[��X   ''r|  G?k�+���X   WRBr}  G?w8N��X   VBZr~  G?�b�O�BX   VBPr  G?��r[��NG?��r[��hMG?�/���X   MDr�  G?���/9X   WPr�  G?r�r[��X   oovr�  G?b�r[��X   RPr�  G?b�r[��X   VBr�  G?k�+���X   JJr�  G?k�+���X   NNPr�  G?k�+���X   ``r�  G?b�r[��uX   WPr�  j  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   DTr�  G?�*⻌ׁX   NNPr�  G?ͼ�<��bX   TOr�  G?�70��#X   VBNr�  G?��� ��X   NNr�  G?��.���X   INr�  G?����|�X   RPr�  G?x��߁�X   PRPr�  G?�C~��nCX   VBGr�  G?�$�E�X   RBr�  G?�|<�]�BX   ``r�  G?n��u� X   PRP$r�  G?p�M�X�X   JJr�  G?�u̡�kX   CCr�  G?SIw�X   CDr�  G?�i���H�X   NNSr�  G?�̡�j��X   JJSr�  G?X��߁�X   VBDr�  G?e��2���X   VBr�  G?o�98�X   VBZr�  G?J�=fڜX   JJRr�  G?^��u� X   oovr�  G?\���3^h�G?>��u� X   RBSr�  G?L���3^X   WRBr�  G?V�X)X   WPr�  G?J�=fڜX   VBPr�  G?6�X)X   ''r�  G?.��u� X   MDr�  G?H��߁�X   NNPSr�  G?T�#�hMG?6�X)X   POSr�  G?6�X)X   WDTr�  G?&�X)uj  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   NNPr�  G?��vsX   JJr�  G?΄R�d�X   NNr�  G?�t�0X   NNSr�  G?���|G�nX   JJSr�  G?�ʵdYI�X   CDr�  G?��` -�X   RBSr�  G?�Ki���X   VBNr�  G?h���[X   oovr�  G?T����X   ``r�  G?s�0���X   INr�  G?m\N�_RX   JJRr�  G?X���[X   VBGr�  G?kY}H�̅X   NNPSr�  G?��W��%X   DTr�  G?d'ja�X   VBr�  G?<�WzxA�X   WDTr�  G?���WX   VBPr�  G?6�l1X   RBr�  G?\'ja�=X   MDr�  G?#N:Q��OX   VBZr�  G?@�lh�G?3N:Q��OX   VBDr�  G?9���WX   WPr�  G?0�lX   CCr�  G?���WX   WRBr�  G?#N:Q��OX   POSr�  G?���WX   TOr�  G?���WX   PRPr�  G?���Wuj�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   POSr�  G?�Uc�a�X   NNPr�  G?���W���X   NNr�  G?ȎO~N��h�G?�M�#�I�X   NNPSr�  G?�pw�rZX   INr�  G?��?�/vX   PRPr�  G?/Ll��rX   CCr�  G?��Vs1{X   NNSr�  G?�����2X   JJr�  G?��,5��X   VBPr�  G?�(����X   VBDr�  G?��R��TX   CDr�  G?�18�+AlX   DTr�  G?]�ͭ�SX   VBNr�  G?��x��zX   JJSr�  G?"�tm�xX   WPr�  G?R�tm�xX   WRBr�  G?E���X   RBr�  G?y�,5��X   TOr�  G?uRv�oA�X   VBGr�  G?`ҭ�-�PX   VBr�  G?��tm�xhMG?����dX   VBZr�  G?�G=����X   ''r�  G?a�$�hX   oovr�  G?fL�B$��NG?E���X   RPr�  G?)	� �X   WDTr�  G?OLl��rX   MDr�  G?a��&��`X   PRP$r�  G?	� �X   JJRr�  G?"�tm�xX   RBSr�  G?"�tm�xX   ``r�  G?Q�$�huX   NNr�  ja  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   VBr�  G?ߚ\���X   NNPr�  G?������'X   VBNr�  G?_E�Z@�h�G?���Z�X   PRP$r�  G?�}��+2/X   DTr   G?�}oC�NX   WDTr  G?z�	<?�X   JJr  G?���S*��X   WPr  G?�؄�7�X   ``r  G?\%U��X   NNSr  G?����5�X   INr  G?���pJFX   PRPr  G?j�	<?�X   WRBr  G?_E�Z@�X   VBGr	  G?�h�[yT}X   NNr
  G?�R�vL�X   RBr  G?�3B6=!X   CDr  G?l%U��X   JJRr  G?I�e��GX   VBDr  G?9�e��GX   NNPSr  G?Y�e��GX   CCr  G?BÎiY�X   TOr  G?BÎiY�X   JJSr  G?9�e��GX   RBSr  G?BÎiY�hMG?BÎiY�NG?OE�Z@�X   oovr  G?BÎiY�uja  j�  �r  h h(h
c__builtin__
__main__
hNN}r  Ntr  Rr  �r  Rr  (h�G?��%o|.X   DTr  G?�`@�8�X   NNPr  G?��"ly+X   PRP$r  G?����vNX   VBNr  G?��X���X   NNr  G?�-sD�-X   WPr   G?������!X   RBr!  G?�4���X   ''r"  G??�(R��X   INr#  G?�6<�qy�X   VBGr$  G?��C!G\�X   JJr%  G?��]�n�X   PRPr&  G?���n0��X   NNSr'  G?�Ex?cX   CDr(  G?{z��5X   RPr)  G?�y�֨zX   ``r*  G?d���+�X   TOr+  G?�Tݍ'�X   CCr,  G?�����^�X   VBr-  G?{z��5X   JJRr.  G?y���$v�X   WRBr/  G?}~e�pX   VBDr0  G?9|��ӫX   JJSr1  G?I|��ӫhMG?o@�+��X   VBPr2  G?9|��ӫX   WDTr3  G?bQ�b�X#X   POSr4  G?3��.��X   oovr5  G?p������X   MDr6  G?3��.��X   RBSr7  G?3��.��NG?Q���@�X   VBZr8  G?I|��ӫX   NNPSr9  G?)|��ӫuj�  h��r:  h h(h
c__builtin__
__main__
hNN}r;  Ntr<  Rr=  �r>  Rr?  (NG?��+ݕ�X   ''r@  G?bҕ:@�h�G?Bҕ:@�X   ``rA  G?_�0�%�X   VBrB  G?Bҕ:@�uX   VBrC  h��rD  h h(h
c__builtin__
__main__
hNN}rE  NtrF  RrG  �rH  RrI  (X   NNPrJ  G?�6b���X   NNrK  G?�ᕋg�h�G?�����X   INrL  G?�d���WX   WPrM  G?������X   DTrN  G?�d���WX   CDrO  G?��ay�\hX   VBGrP  G?�H��2X   RBrQ  G?v���DX   JJrR  G?��+E��X   NNSrS  G?�N<S"�X   PRP$rT  G?��MjbX   WRBrU  G?p8Ʒ�G�X   WDTrV  G?k���ċX   JJRrW  G?r��'-�X   PRPrX  G?�%p���X   TOrY  G?v���DX   VBNrZ  G?k���ċhMG?b��'-�X   VBr[  G?W,��p�X   ''r\  G?B��'-�X   NNPSr]  G?R��'-�X   ``r^  G?b��'-�X   JJSr_  G?`8Ʒ�G�X   VBZr`  G?B��'-�X   CCra  G?W,��p�X   MDrb  G?B��'-�X   oovrc  G?b��'-�NG?B��'-�X   VBDrd  G?B��'-�uh�jJ  �re  h h(h
c__builtin__
__main__
hNN}rf  Ntrg  Rrh  �ri  Rrj  (X   POSrk  G?��B~Vq
h�G?���۲�hMG?���ʠX   VBPrl  G?��H��X   RBrm  G?{~�v�,MX   NNPrn  G?�$MF�|sX   CDro  G?��hR��X   CCrp  G?��p���X   ''rq  G?d �&^YQX   NNPSrr  G?hp�����X   VBDrs  G?�"�:�GX   INrt  G?���c�X   NNru  G?��W���X   VBGrv  G?p,��X   MDrw  G?o��X   VBZrx  G?��:h�{X   TOry  G?�C�`%aPX   JJrz  G?vHȏuX   NNSr{  G?����{�X   VBr|  G?{P�ؤ��X   PRPr}  G?T �&^YQX   WDTr~  G?j<�$MF�X   WRBr  G?Z��`jc�X   VBNr�  G?|���X   oovr�  G?l���NG?kP�ؤ��X   DTr�  G?d|�b{vWX   WPr�  G?T �&^YQX   PRP$r�  G?' �GA�X   RBSr�  G?' �GA�X   ``r�  G?A@�Euq!X   JJSr�  G?,���X   JJRr�  G? �GA�uX   NNPr�  h��r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (NG?��첉LX   NNr�  G?Qӄ��X   ''r�  G?]�&��(X   CDr�  G?`��� �X   WPr�  G?#t_r�K�X   NNPr�  G?i�C�eSX   VBDr�  G?)�C�eSX   ``r�  G?A�W~�E�X   oovr�  G?)�C�eSX   INr�  G?6�o[rX�h�G?N͗ �xSX   VBNr�  G?�C�eSX   CCr�  G?)�C�eSX   VBr�  G?)�C�eSX   NNSr�  G?#t_r�K�X   VBZr�  G?�C�eSX   DTr�  G?�C�eShMG?#t_r�K�X   POSr�  G?�C�eSX   VBGr�  G?�C�eSuX   NNr�  j  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   VBDr�  G?��)��X   INr�  G?��Kz�NX   NNPr�  G?̀ʰLX   POSr�  G?�5��0��X   NNr�  G?�I^{�nQX   ''r�  G?u���h�G?�;+HPX   VBZr�  G?��h��1X   CCr�  G?���R޿X   TOr�  G?�\�"�MX   JJr�  G?m��(X   VBNr�  G?�yf톙X   MDr�  G?s � 2�X   WDTr�  G?e���X   RBr�  G?��Kz�NX   VBr�  G?�ǅ��X   NNSr�  G?��U�`hMG?�dI囶X   NNPSr�  G?m��(X   CDr�  G?w9���DX   VBGr�  G?s � 2�X   oovr�  G?`�U�`X   VBPr�  G?�9���DX   DTr�  G?}��(X   WRBr�  G?e���NG?m��(X   PRPr�  G?iV	�C�X   ``r�  G?`�U�`X   RBSr�  G?P�U�`uj  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   INr�  G?Ƅ��ڕX   TOr�  G?��t��vh�G?�L����rX   DTr�  G?��#�ُiX   VBNr�  G?�;�<<�aX   PRP$r�  G?�"� �5jX   WPr�  G?���J�1X   RBr�  G?���`y�X   VBDr�  G?`��]��3X   WDTr�  G?�T����X   WRBr�  G?~S�p�S6X   NNr�  G?��庠Z�X   CDr�  G?t�^��bX   NNSr�  G?�<�CI�X   NNPr�  G?�["'��gX   RPr�  G?�C�B�X   JJr�  G?�&6\��X   JJSr�  G?]:W��{X   VBGr�  G?�+��`��X   VBr�  G?q���=}X   JJRr�  G?U����oX   oovr�  G?e����oX   PRPr�  G?�͋8�X   CCr�  G?hC�B�hMG?m:W��{X   MDr�  G?=:W��{X   NNPSr�  G?HC�B�X   ''r�  G?3hя���X   ``r�  G?Z� %�X   VBZr�  G?HC�B�X   RBSr�  G?Chя���NG?HC�B�uj�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   DTr�  G?�2\S�6�X   PRP$r�  G?��o�`4X   WPr�  G?�����X   NNPr�  G?�D�"��X   PRPr�  G?�R*�ɩ�X   WDTr�  G?���F��h�G?�����X   VBNr�  G?\E�Pf}X   INr�  G?�����X   CDr�  G?�`�K�}�X   VBGr�  G?�Ե$�X   WRBr�  G?v��SE�X   JJr�  G?�o�wFX   TOr�  G?tR*�ɩ�X   VBDr�  G?q���@#X   NNr�  G?�w���X   JJSr�  G?a���@#X   ``r�  G?o΅�sL�X   NNSr�  G?�B���X   RBr�  G?|E�Pf}X   oovr�  G?q���@#hMG?Q���@#X   JJRr�  G?e4Y<L��X   MDr   G?<E�Pf}X   NNPSr  G?X��Y�dX   VBZr  G?Q���@#X   CCr  G?E4Y<L��NG?U4Y<L��X   VBr  G?E4Y<L��X   VBPr  G?<E�Pf}uj�  j�  �r  h h(h
c__builtin__
__main__
hNN}r  Ntr  Rr	  �r
  Rr  (X   NNr  G?��~3���X   RBSr  G?nhb� |�X   DTr  G?W�_�0,X   CDr  G?��"�i��X   NNSr  G?��6DhsX   JJr  G?�J��GX   NNPr  G?���ֹ-�X   VBGr  G?t[���mX   JJSr  G?�8�#k
X   ``r  G?n��{3�X   INr  G?l�a� 2�X   RBr  G?_��f�X   JJRr  G?b�>�X   NNPSr  G?)b�p��X   PRP$r  G?$�vY.rh�G?M&�k��X   VBNr  G?k��º��X   WPr  G?S]�nR�X   WDTr  G?( 
��"X   oovr  G?K$��1�X   VBZr  G?4�vY.rX   PRPr   G?0\^���X   POSr!  G? 
��"X   TOr"  G?$�vY.rX   MDr#  G?4�vY.rX   VBDr$  G?@\^���X   VBPr%  G?( 
��"hMG?\^���X   CCr&  G?\^���NG?\^���ujb  j�  �r'  h h(h
c__builtin__
__main__
hNN}r(  Ntr)  Rr*  �r+  Rr,  (X   NNPr-  G?ڋ��h��X   DTr.  G?�]lPD�qX   PRP$r/  G?�챶(:X   WPr0  G?�E>�VL0X   WDTr1  G?qm�r��X   CDr2  G?�,�F	qh�G?��#)�X   JJSr3  G?Uo����X   VBGr4  G?��C��X   ``r5  G?iUǪ~~!X   NNr6  G?���2҉X   INr7  G?��<�?�-X   VBDr8  G?Uo����X   JJr9  G?��ɼ��$X   NNSr:  G?�\S��e�X   RBr;  G?h\S��e�X   PRPr<  G?������SX   NNPSr=  G?};��V�MX   WRBr>  G?`����=X   VBNr?  G?[H���7X   CCr@  G?C}�9��X   oovrA  G?`����=X   TOrB  G?_.��cX   VBZrC  G?Gb߱M
X   VBPrD  G?/.��chMG?7b߱M
NG?7b߱M
X   JJRrE  G??.��cX   MDrF  G?/.��cuX   WRBrG  h>�rH  h h(h
c__builtin__
__main__
hNN}rI  NtrJ  RrK  �rL  RrM  (X   NNPrN  G?�\J���X   VBDrO  G?�f��k/X   NNSrP  G?�V�
�X   INrQ  G?�q��PjX   VBZrR  G?��~��X   JJrS  G?�����KX   NNrT  G?�C[�'X   JJRrU  G?u��&1�6X   VBNrV  G?s��rQ�X   DTrW  G?f8�ꓴX   VBGrX  G?V8�ꓴX   MDrY  G?w�c��/X   VBPrZ  G?��0L�yX   TOr[  G?Xq���խh�G?pU"��IX   NNPSr\  G?���%8�X   CDr]  G?hq���խX   ``r^  G?Xq���խX   RBr_  G?�8��h�EX   oovr`  G?O:x{��X   PRPra  G?O:x{��X   VBrb  G?J�{B��NG?1���"�X   JJSrc  G?1���"�X   WRBrd  G?1���"�hMG?:�{B��X   PRP$re  G?1���"�X   CCrf  G?A���"�uh>jN  �rg  h h(h
c__builtin__
__main__
hNN}rh  Ntri  Rrj  �rk  Rrl  (X   NNSrm  G?�
��{~X   NNPrn  G?ɮ�,��/X   ''ro  G?r\ �!b�h�G?Ŏs��X   NNrp  G?�P���X   INrq  G?�$,^�	fX   VBDrr  G?����˧X   NNPSrs  G?��L��`X   VBZrt  G?�y\f�`�X   POSru  G?�Þ��<X   VBPrv  G?�Ht�aQX   CCrw  G?��~�6�|X   MDrx  G?q|O�+��X   TOry  G?��4��b#X   VBNrz  G?���җ�X   JJr{  G?��{��X   WPr|  G?_y\f�`�X   RBr}  G?�����X   DTr~  G?t�%/nX   VBr  G?��~�6�|X   oovr�  G?d�����NG?T�����X   WDTr�  G?a|O�+��X   WRBr�  G?D�����X   VBGr�  G?a|O�+��hMG?�
��{~X   ``r�  G?[�>�ǎX   CDr�  G?v�4��b#X   PRPr�  G?K�>�ǎX   PRP$r�  G?;�>�ǎujN  jm  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   VBDr�  G?���G|tX   VBZr�  G?�OFr��XX   INr�  G?��:T�fxX   NNr�  G?�X��a˺X   VBPr�  G?��R�[d8h�G?��e��]X   RBr�  G?��ۦ��`X   CCr�  G?���JX   VBr�  G?���a{�X   RPr�  G?P�ۦ��`X   NNPr�  G?�X   VBGr�  G?��1T�X   WDTr�  G?�;�����hMG?�
6Y��X   JJr�  G?�c�k��X   JJRr�  G?V'ψ��X   MDr�  G?�X   TOr�  G?��0J�\nX   VBNr�  G?��z��+rX   NNSr�  G?~v�\A�0X   WPr�  G?w�L�x��X   RBSr�  G?P�ۦ��`X   ''r�  G?[��k$��X   DTr�  G?}@c�%�X   PRP$r�  G?P�ۦ��`X   WRBr�  G?`�ۦ��`X   POSr�  G?��ۦ��`X   oovr�  G?cb՗���X   CDr�  G?P�ۦ��`NG?h��zEX   PRPr�  G?F'ψ��uX   INr�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   JJr�  G?ʂ�A�X   NNr�  G?�Jm1�|X   CDr�  G?��\5bF_X   INr�  G?ci���HX   NNSr�  G?Ġ&��X   NNPr�  G?��ǴJ�X   JJRr�  G?WKw$��X   RBr�  G?ci���HX   JJSr�  G?�-`Uj
1X   VBGr�  G?wKw$��X   VBDr�  G?_I�0�X   MDr�  G?WKw$��X   RBSr�  G?OI�0�X   WPr�  G?ci���HX   VBNr�  G?uZ��AX   CCr�  G?ci���HX   VBZr�  G?WKw$��hMG?OI�0�X   ``r�  G?gKw$��X   DTr�  G?OI�0�X   POSr�  G?WKw$��uj�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   NNr�  G?㒐�U�X   NNPr�  G?��g��X   ``r�  G?oDe�JBqX   VBr�  G?oDe�JBqX   JJr�  G?�����i�hMG?_De�JBqX   NNSr�  G?Ʒ���FX   RBr�  G?oDe�JBqX   CDr�  G?��U�sLX   VBNr�  G?{[���#X   INr�  G?��y)	�`X   WPr�  G?{[���#h�G?���U�sX   CCr�  G?s����i�X   VBGr�  G?s����i�X   VBZr�  G?_De�JBqX   JJSr�  G?_De�JBqX   NNPSr�  G?oDe�JBqX   TOr�  G?gsL6���X   RPr�  G?_De�JBqX   DTr�  G?_De�JBqX   MDr�  G?_De�JBquh{jL  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   INr�  G?ť}�$h�G?�u�Z
X   NNr�  G?�НSրX   VBDr�  G?����.�|X   JJr�  G?�d�m=��X   POSr�  G?��E���X   CCr�  G?�T,���5X   ``r�  G?p&���tX   VBNr�  G?�����sX   NNPr�  G?�HX�lhMG?�C���o�X   NNSr�  G?�E����*X   VBr�  G?�&���tX   RBr�  G?�)7�hN�X   VBZr�  G?����N:�X   TOr�  G?��7vE4X   WPr�  G?j��m�!X   PRPr�  G?L�^S�X   WDTr�  G?r׭�J\X   WRBr�  G?i���c&X   VBPr�  G?�&���tX   VBGr�  G?|�^S�X   DTr�  G?q����kdX   MDr�  G?t�˼MX   CDr�  G?\�^S�X   RBSr�  G?L�^S�X   ''r�  G?`&���tX   oovr�  G?U�ƾT�ENG?L�^S�X   PRP$r�  G?<�^S�uX   POSr   jM  �r  h h(h
c__builtin__
__main__
hNN}r  Ntr  Rr  �r  Rr  (X   NNr  G?����X   VBGr  G?c�*�`X   JJr	  G?�(c�Z�X   NNSr
  G?�U��rh�G?�	��bX   PRPr  G?S�*�`hMG?p��%k�X   VBNr  G?�ѫ��:X   CCr  G?w�:5u�X   VBr  G?S�*�`X   NNPr  G?���|#�WX   RBSr  G?l��@&�X   INr  G?s�*�`X   NNPSr  G?g�:5u�X   ``r  G?\��@&�X   CDr  G?ub0��X   RBr  G?g�:5u�X   DTr  G?S�*�`X   JJSr  G?w�:5u�X   VBPr  G?\��@&�X   TOr  G?\��@&�X   VBDr  G?\��@&�X   oovr  G?S�*�`X   VBZr  G?S�*�`uX   NNr  hM�r  h h(h
c__builtin__
__main__
hNN}r  Ntr   Rr!  �r"  Rr#  (X   WPr$  G?�(���"X   INr%  G?���e�X�X   VBDr&  G?����)5oX   ``r'  G?���q�)X   VBGr(  G?��1��X   NNPr)  G?�ಿ.�dX   VBNr*  G?���q�)X   CDr+  G?j���A�X   RBr,  G?�s�����X   WRBr-  G?���0-7X   DTr.  G?��x��\X   NNr/  G?�tƏ��]X   JJr0  G?���q�)X   CCr1  G?��a� 
X   WDTr2  G?�K[*C=�X   NNSr3  G?��}��hX   PRP$r4  G?T<H�1SX   VBZr5  G?�#3����X   VBPr6  G?���q�)X   PRPr7  G?�#3����X   VBr8  G?j���A�X   oovr9  G?|���]E�X   MDr:  G?z���A�X   JJRr;  G?g��k�9�X   ''r<  G?d<H�1SX   TOr=  G?g��k�9�X   JJSr>  G?J���A�hMG?J���A�NG?J���A�h�G?J���A�uhMj$  �r?  h h(h
c__builtin__
__main__
hNN}r@  NtrA  RrB  �rC  RrD  (X   JJrE  G?�(����X   VBPrF  G?���+/�X   VBDrG  G?вB�YX   CDrH  G?x����X   RBrI  G?�����X   NNrJ  G?�U{SArlX   VBZrK  G?˶��8�X   NNPrL  G?�^��\��X   MDrM  G?�����X   NNSrN  G?�����X   INrO  G?\~q�ΕX   VBrP  G?h����X   VBGrQ  G?h����X   DTrR  G?U^��\��X   PRPrS  G?U^��\��X   WPrT  G?U^��\��h�G?U^��\��X   ``rU  G?L~q�ΕX   WRBrV  G?L~q�ΕX   JJRrW  G?L~q�Εuj$  jE  �rX  h h(h
c__builtin__
__main__
hNN}rY  NtrZ  Rr[  �r\  Rr]  (X   NNr^  G?���9��$X   NNSr_  G?�yq[���X   NNPr`  G?�N���OX   VBDra  G?����n�X   JJrb  G?�W�4�X   VBGrc  G?�EX5-X   CDrd  G?iޕ��j�X   VBZre  G?���'��X   TOrf  G?V���	�X   VBPrg  G?V���	�X   RBrh  G?V���	�X   CCri  G?a?�4G$X   MDrj  G?F���	�X   VBNrk  G?\�m���hMG?Q?�4G$h�G?o�EX5-X   INrl  G?\�m���X   ``rm  G?F���	�X   NNPSrn  G?F���	�X   DTro  G?F���	�X   JJRrp  G?F���	�uNh�rq  h h(h
c__builtin__
__main__
hNN}rr  Ntrs  Rrt  �ru  Rrv  (X   NNrw  G?�
��%~X   JJSrx  G?C���ܼX   NNPry  G?�I�~5�DX   JJrz  G?��AZD�X   CDr{  G?�s�jɊ?X   INr|  G?�ۗm� X   NNSr}  G?�6'�t�X   TOr~  G?�k�O�hX   VBZr  G?����3}X   VBGr�  G?y��m9��X   VBDr�  G?q�H�$X   NNPSr�  G?e�9�SX   CCr�  G?m?��fKhMG?S���ܼX   RBr�  G?c���ܼX   VBNr�  G?M?��fKX   JJRr�  G?]?��fKX   VBPr�  G?c���ܼX   WPr�  G?C���ܼuNh �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   VBr�  G?�������X   WPr�  G?�H����X   WDTr�  G?�X�~��zX   DTr�  G?�	K1�"�X   WRBr�  G?�	K1�"�X   NNPr�  G?{	K1�"�X   RBr�  G?{	K1�"�uX   NNPr�  hM�r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   WRBr�  G?� mh�5lX   VBDr�  G?�9D����X   NNPr�  G?�߄�4#�X   WDTr�  G?�\PX�X   NNSr�  G?��-�ýTX   VBNr�  G?��Џ�m�X   INr�  G?��磯�X   NNr�  G?�֋SV�X   VBr�  G?t���FX   CDr�  G?���x�W�X   WPr�  G?Жo�)t�X   CCr�  G?�d܇@X   DTr�  G?� mh�5lX   VBZr�  G?�4����`X   PRP$r�  G?T���FX   JJSr�  G?T���FX   RBr�  G?�^sdoXX   VBGr�  G?�9D��X   JJr�  G?�[��/�X   MDr�  G?r��%.��X   ``r�  G?n�r�i#X   NNPSr�  G?T���FX   TOr�  G?v9D����X   VBPr�  G?kZ-M[X   oovr�  G?d���FX   ''r�  G?a\PX�X   PRPr�  G?q\PX�h�G?d���FNG?KZ-M[uhMj�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   JJr�  G?�ص��D�X   VBDr�  G?��Ȕ�X   VBNr�  G?����&vHX   MDr�  G?�U2
��HX   RBr�  G?�:P;���X   VBZr�  G?���D=5X   VBPr�  G?��p}��lX   INr�  G?����&vHX   DTr�  G?�w�u
V�X   VBr�  G?s����#X   CCr�  G?jw�u
V�X   PRPr�  G?�(�i�X   VBGr�  G?zw�u
V�X   NNPr�  G?jw�u
V�X   NNSr�  G?jw�u
V�X   PRP$r�  G?jw�u
V�uj�  jO  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   NNPr�  G?�rkx.X   ``r�  G?jWAh�JX   DTr�  G?јHo��_X   PRPr�  G?�WAh�JX   NNr�  G?�+���EX   INr�  G?�)��ΜX   CDr�  G?��pŎg�X   VBNr�  G?��o WAX   NNSr�  G?�t�0���X   TOr�  G?�v���VnX   VBGr�  G?�v���VnX   RBr�  G?�v���VnX   JJr�  G?�����X   VBr�  G?zWAh�JX   PRP$r�  G?�v���VnX   WPr�  G?�v���Vnh�G?s�pŎg�X   WDTr�  G?jWAh�JX   RPr�  G?jWAh�JX   VBDr�  G?s�pŎg�X   JJSr�  G?s�pŎg�NG?jWAh�JX   WRBr�  G?jWAh�JX   oovr�  G?s�pŎg�X   VBZr�  G?jWAh�JhMG?jWAh�JuX   VBr�  h��r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   JJr�  G?�+�Djz�X   NNr�  G?�Ʉ�i�X   CDr�  G?��%QZOh�G?g�%QZOX   NNSr�  G?�%�
���X   NNPr�  G?��]�)LX   ``r�  G?{�+���X   JJSr�  G?�ڮ����X   RBr�  G?g�%QZOX   VBGr�  G?��%QZOX   INr�  G?g�%QZOX   RBSr�  G?g�%QZOX   VBNr�  G?o�1�;�X   JJRr�  G?_�1�;�X   MDr�  G?_�1�;�uj�  jn  �r 	  h h(h
c__builtin__
__main__
hNN}r	  Ntr	  Rr	  �r	  Rr	  (X   NNr	  G?���~�UhMG?�T��uh�G?ͼ� ���X   NNPr	  G?��ŧ��X   INr	  G?����-mX   DTr		  G?�6J��(�X   CCr
	  G?���1{\oX   PRPr	  G?f���ɀX   POSr	  G?�7po0X   CDr	  G?r���HX   ''r	  G?r���HX   TOr	  G?�c+���{X   VBNr	  G?�N �X   VBPr	  G?��k��r�X   VBDr	  G?��	��lX   VBZr	  G?��mz�PX   VBr	  G?�\�*��X   VBGr	  G?q��Z��X   WDTr	  G?YJmҁ�X   WRBr	  G?b$���_uX   WPr	  G?R$���_uX   NNSr	  G?�+�P��X   JJr	  G?~��t�tX   MDr	  G?d�p���X   RBr	  G?���t�tX   ``r	  G?a3���	NG?Z���X   RBSr	  G?%��1{\oX   NNPSr	  G?U��1{\oX   oovr 	  G?i�-mWYiX   JJSr!	  G?E��1{\oX   JJRr"	  G?%��1{\oX   PRP$r#	  G?%��1{\ouX   PRP$r$	  j�  �r%	  h h(h
c__builtin__
__main__
hNN}r&	  Ntr'	  Rr(	  �r)	  Rr*	  (X   CCr+	  G?���f���h�G?׌3H_��X   NNr,	  G?��6-~hMG?���p�X   INr-	  G?�      X   TOr.	  G?���f���X   DTr/	  G?w(�i�X   ``r0	  G?s����#X   RBr1	  G?�4nlX   VBDr2	  G?��RL��X   WPr3	  G?c����#X   POSr4	  G?���f���X   NNPr5	  G?�4nlX   WRBr6	  G?jw�u
V�X   VBNr7	  G?���p�X   VBGr8	  G?nlZ�G"X   NNSr9	  G?�1���scX   VBZr:	  G?��-�N�X   MDr;	  G?x�p}��lX   CDr<	  G?S����#X   VBPr=	  G?`���&vHX   VBr>	  G?x�p}��lX   RPr?	  G?S����#X   ''r@	  G?S����#X   JJrA	  G?c����#X   oovrB	  G?Jw�u
V�NG?Zw�u
V�X   WDTrC	  G?`���&vHX   PRPrD	  G?Jw�u
V�uj�  j�  �rE	  h h(h
c__builtin__
__main__
hNN}rF	  NtrG	  RrH	  �rI	  RrJ	  (X   INrK	  G?�V��0.X   DTrL	  G?��ݦ�@X   CDrM	  G?bq0K�ߜh�G?�=Q��6X   TOrN	  G?�2�H��*X   NNrO	  G?��VU{�X   CCrP	  G?�Ѫu9X   NNSrQ	  G?��iY�I�X   RBrR	  G?���:pD<X   NNPrS	  G?tIN����X   VBNrT	  G?�q0K�ߜX   VBPrU	  G?rq0K�ߜX   VBrV	  G?�ZMW|$X   JJRrW	  G?p�ݦ�@hMG?���:pD<X   VBGrX	  G?���z-�X   ''rY	  G?f!m'�UX   POSrZ	  G?v!m'�UX   VBDr[	  G?w���"�X   VBZr\	  G?yѪu9X   WRBr]	  G?p�ݦ�@X   JJr^	  G?v!m'�UX   WPr_	  G?]���ae�X   MDr`	  G?m���ae�X   WDTra	  G?iѪu9X   oovrb	  G?V!m'�UNG?bq0K�ߜX   PRPrc	  G?bq0K�ߜX   PRP$rd	  G?M���ae�X   ``re	  G?V!m'�UuX   VBDrf	  j�  �rg	  h h(h
c__builtin__
__main__
hNN}rh	  Ntri	  Rrj	  �rk	  Rrl	  (X   INrm	  G?֜�OF�X   VBDrn	  G?�֓8�XX   NNro	  G?��\���{h�G?��~��X   WRBrp	  G?��{as�X   VBZrq	  G?���\�X   TOrr	  G?�Oޟ$�X   NNPrs	  G?��m��EpX   NNSrt	  G?���q?zX   VBru	  G?��{as�X   VBNrv	  G?�#�4'V�X   POSrw	  G?�9���gX   CDrx	  G?��\�<�X   VBGry	  G?�uJ͢lX   MDrz	  G?l�)�-�X   RBr{	  G?��K����X   JJr|	  G?s�{as�X   CCr}	  G?�I��QX   WDTr~	  G?s�{as�hMG?�uJ͢lX   VBPr	  G?c�{as�X   WPr�	  G?g�x9��X   DTr�	  G?p�m��EpX   PRP$r�	  G?S�{as�X   RBSr�	  G?c�{as�X   ``r�	  G?\�)�-�X   PRPr�	  G?S�{as�ujm	  j�  �r�	  h h(h
c__builtin__
__main__
hNN}r�	  Ntr�	  Rr�	  �r�	  Rr�	  (X   INr�	  G?�6�%���X   VBDr�	  G?�
Ji��X   CDr�	  G?�-��h�G?�9��6X   TOr�	  G?�	ܥ2M�X   VBZr�	  G?�q�(C�X   CCr�	  G?�����X   NNSr�	  G?��(���X   NNr�	  G?��h'r��X   VBNr�	  G?�ט����hMG?��w\ԙX   VBGr�	  G?u4|�fHwX   POSr�	  G?tD���.�X   NNPr�	  G?~�dX   DTr�	  G?l��-�X   PRPr�	  G?M��c9 X   VBPr�	  G?�s��j�X   WDTr�	  G?|`���&X   MDr�	  G?�w���;X   WRBr�	  G?i�����X   JJr�	  G?z���ڔX   RBr�	  G?�-��X   VBr�	  G?Z1�����X   WPr�	  G?]��c9 X   ''r�	  G?rf���X   oovr�	  G?X�tZү�X   ``r�	  G?Fs��j�X   JJRr�	  G?3�)�B&NG?av����SX   RPr�	  G?#�)�B&X   RBSr�	  G?#�)�B&X   JJSr�	  G?#�)�B&X   PRP$r�	  G?#�)�B&X   NNPSr�	  G?#�)�B&uX   NNr�	  j�  �r�	  h h(h
c__builtin__
__main__
hNN}r�	  Ntr�	  Rr�	  �r�	  Rr�	  (X   NNPr�	  G?�㪀?��X   VBNr�	  G?��(C��X   INr�	  G?�R�9���X   DTr�	  G?ş��w�X   NNr�	  G?��W��X   VBDr�	  G?��(C��X   TOr�	  G?�!�L�X   WPr�	  G?��16.��X   JJr�	  G?��j`oYX   NNSr�	  G?��	�^rh�G?�\��&F�X   WRBr�	  G?o�G��jX   PRP$r�	  G?��:(�۶X   PRPr�	  G?�����X   RPr�	  G?��(C��X   RBr�	  G?���W��X   MDr�	  G?_�G��jX   JJRr�	  G?o�G��jX   NNPSr�	  G?_�G��jX   CDr�	  G?w�5�x��X   VBGr�	  G?g�5�x��X   VBZr�	  G?w�5�x��X   WDTr�	  G?o�G��jNG?_�G��jX   ``r�	  G?s�,��X   CCr�	  G?g�5�x��X   JJSr�	  G?_�G��jX   oovr�	  G?g�5�x��X   ''r�	  G?g�5�x��X   VBr�	  G?g�5�x��hMG?_�G��juj�  j�	  �r�	  h h(h
c__builtin__
__main__
hNN}r�	  Ntr�	  Rr�	  �r�	  Rr�	  (X   NNPr�	  G?˟׃)��X   POSr�	  G?�]��rKhMG?�ޮ�[��X   VBNr�	  G?�ޮ�[��h�G?��5#�3X   NNSr�	  G?���l��X   INr�	  G?�v�8��X   NNr�	  G?�>k��aX   TOr�	  G?��'���X   VBDr�	  G?������X   CCr�	  G?�]��rKX   oovr�	  G?���*,��X   VBGr�	  G?�ޮ�[��X   RBr�	  G?���*,��X   VBZr�	  G?z��*,��X   VBPr�	  G?z��*,��X   MDr�	  G?t>k��aX   JJRr�	  G?j��*,��X   CDr�	  G?�>k��aX   PRPr�	  G?j��*,��X   JJr�	  G?��'���NG?j��*,��X   DTr�	  G?t>k��aX   VBr�	  G?t>k��aX   ``r�	  G?j��*,��uhMj�  �r�	  h h(h
c__builtin__
__main__
hNN}r�	  Ntr�	  Rr�	  �r�	  Rr�	  (X   NNPr�	  G?�A}��X   VBNr�	  G?�SYMe5�X   WRBr�	  G?��Gq�wX   WDTr�	  G?��_A}�X   DTr�	  G?�Gq�wX   NNr�	  G?�_A}�X   TOr�	  G?��w�GqX   RBr�	  G?��_A}�X   INr�	  G?��_A}�X   NNSr�	  G?��_A}�X   JJr�	  G?��Gq�wX   RPr�	  G?��_A}�X   WPr�	  G?��SYMe6X   CCr�	  G?��Gq�whMG?��Gq�wX   VBGr�	  G?��_A}�h�G?��_A}�X   PRPr�	  G?��SYMe6X   PRP$r 
  G?��Gq�wX   VBZr
  G?��_A}�X   CDr
  G?��_A}�X   JJSr
  G?��_A}�uX   NNPr
  jn  �r
  h h(h
c__builtin__
__main__
hNN}r
  Ntr
  Rr
  �r	
  Rr

  (X   PRP$r
  G?�M�h��X   NNPr
  G?�1^'���h�G?����薦X   INr
  G?�o��[�X   VBNr
  G?��&�D�X   VBr
  G?pII�d�X   DTr
  G?�1^'���X   WPr
  G?�r�N��uX   VBZr
  G?|�A%'0ZX   TOr
  G?�:�a5pzX   JJr
  G?��c��X   NNSr
  G?��A�qX   VBDr
  G?vd�x�ʐX   VBGr
  G?��A%'0ZX   WDTr
  G?d[�?��X   NNr
  G?�5��t
.X   RBr
  G?��,Ɋ�>X   PRPr
  G?��{*>iX   oovr
  G?|�A%'0ZX   MDr
  G?d[�?��X   RPr
  G?�m�!�(X   RBSr
  G?Xm�!�(X   JJRr 
  G?pII�d�X   CDr!
  G?�r�N��uX   WRBr"
  G?rRs�1^X   ``r#
  G?d[�?��X   JJSr$
  G?rRs�1^X   CCr%
  G?Xm�!�(hMG?PII�d�NG?`II�d�X   VBPr&
  G?Xm�!�(X   POSr'
  G?Xm�!�(X   ''r(
  G?PII�d�ujn  j
  �r)
  h h(h
c__builtin__
__main__
hNN}r*
  Ntr+
  Rr,
  �r-
  Rr.
  (X   NNr/
  G?�������X   NNSr0
  G?ОZ�	�X   VBNr1
  G?��}�pX   JJr2
  G?�&��A�jX   JJSr3
  G?���0�X�X   DTr4
  G?|�m���X   CDr5
  G?��m���X   NNPr6
  G?��}�puX   JJr7
  j  �r8
  h h(h
c__builtin__
__main__
hNN}r9
  Ntr:
  Rr;
  �r<
  Rr=
  (X   NNr>
  G?Ҕ�)JR�X   NNSr?
  G?�fٶm�gh�G?�� HX   NNPr@
  G?���xX   TOrA
  G?��!B�X   VBNrB
  G?��!�r�X   JJrC
  G?���xX   DTrD
  G?���xX   INrE
  G?�� HX   VBDrF
  G?�� HX   ''rG
  G?��`X   VBZrH
  G?��`X   VBrI
  G?�� HX   ``rJ
  G?�� HX   PRPrK
  G?�� HX   RBrL
  G?��`X   WPrM
  G?�� HX   oovrN
  G?x�`X   CCrO
  G?x�`X   VBPrP
  G?x�`X   CDrQ
  G?x�`uj  j>
  �rR
  h h(h
c__builtin__
__main__
hNN}rS
  NtrT
  RrU
  �rV
  RrW
  (hMG?���7^�h�G?���W'�DX   ''rX
  G?���W'�DX   RBrY
  G?�g�d$��X   VBDrZ
  G?���7^�X   INr[
  G?��6���{X   CCr\
  G?�=�#4K2X   VBZr]
  G?�ne�g8eX   NNr^
  G?�ckR_X   NNPr_
  G?{W��=��X   NNSr`
  G?�{b��՞X   TOra
  G?�{b��՞X   JJrb
  G?�W��=��X   VBNrc
  G?�g�d$��X   VBGrd
  G?���=.$;X   DTre
  G?pg�d$��X   JJRrf
  G?`g�d$��X   MDrg
  G?���W'�DX   VBrh
  G?e��017�X   oovri
  G?e��017�X   VBPrj
  G?{W��=��NG?`g�d$��X   JJSrk
  G?U��017�X   WDTrl
  G?~��C��X   POSrm
  G?{W��=��X   WPrn
  G?U��017�X   RPro
  G?`g�d$��X   WRBrp
  G?kW��=��X   PRP$rq
  G?U��017�X   RBSrr
  G?U��017�X   PRPrs
  G?U��017�X   ``rt
  G?U��017�X   CDru
  G?U��017�uhMj%  �rv
  h h(h
c__builtin__
__main__
hNN}rw
  Ntrx
  Rry
  �rz
  Rr{
  (X   CDr|
  G?��2��kX   WDTr}
  G?�6zt���X   NNPr~
  G?���z�X   oovr
  G?�$(F޼X   DTr�
  G?ű��Rp�X   NNr�
  G?���/��X   INr�
  G?��ੳӥX   WPr�
  G?ƨ���mX   WRBr�
  G?�-Qy�@X   PRPr�
  G?����}Y1X   PRP$r�
  G?�$(F޼X   NNSr�
  G?��ੳӥX   VBNr�
  G?����}Y1X   JJSr�
  G?�$(F޼X   VBGr�
  G?�[_u'X   JJr�
  G?�H�jdGX   RBr�
  G?�H�jdGh�G?n�ੳӥX   JJRr�
  G?n�ੳӥX   TOr�
  G?n�ੳӥX   MDr�
  G?n�ੳӥuj%  j|
  �r�
  h h(h
c__builtin__
__main__
hNN}r�
  Ntr�
  Rr�
  �r�
  Rr�
  (h�G?�p�|�3X   NNSr�
  G?�������hMG?��2�o?X   INr�
  G?����X   TOr�
  G?��h�d�X   JJr�
  G?��m���X   VBNr�
  G?Uq�<Pk:X   NNr�
  G?��(5��X   NNPr�
  G?�0@UǴ�X   WPr�
  G?�sD[$0@X   VBDr�
  G?��-� +X   CDr�
  G?ql��WX   WDTr�
  G?��W��X   CCr�
  G?�����#X   WRBr�
  G?z"�!��X   JJRr�
  G?5q�<Pk:NG?�%�_)�X   ``r�
  G?@q�<PkX   VBZr�
  G?d�h�d�X   POSr�
  G?r *��yX   DTr�
  G?ywI��TX   VBPr�
  G?Rï��]�X   VBGr�
  G?f�q�X   RBr�
  G?]|�2�oX   NNPSr�
  G?@q�<PkX   oovr�
  G?Z�h�d�X   MDr�
  G?Rï��]�X   VBr�
  G?Pq�<PkX   JJSr�
  G?Eq�<Pk:X   PRPr�
  G?J�h�d�uj|
  h��r�
  h h(h
c__builtin__
__main__
hNN}r�
  Ntr�
  Rr�
  �r�
  Rr�
  (NG?��䎊q�X   ''r�
  G?J6��C-h�G?J6��C-uX   WPr�
  j  �r�
  h h(h
c__builtin__
__main__
hNN}r�
  Ntr�
  Rr�
  �r�
  Rr�
  (X   NNPr�
  G?�2�m���X   DTr�
  G?✗�3�SX   VBNr�
  G?�g�'�@X   NNr�
  G?�	
KZ>�X   PRPr�
  G?�K�m�`XX   VBDr�
  G?���}�X   INr�
  G?���d|�JX   JJr�
  G?�K�m�`XX   VBPr�
  G?��|�4��X   VBr�
  G?��ƒ6BX   TOr�
  G?����GX   VBGr�
  G?��d��O�X   MDr�
  G?[ޠI�mX   WPr�
  G?6K�m�`XX   JJRr�
  G?\��L��X   RBr�
  G?���{W.X   RPr�
  G?a�)$}�X   CDr�
  G?��g��\X   WRBr�
  G?kޠI�mX   NNSr�
  G?��r�X   ``r�
  G?t���1��X   oovr�
  G?Y��$t��X   VBZr�
  G?{�[Nѝh�G?FK�m�`XX   PRP$r�
  G?U.P�U��X   JJSr�
  G?J�=���X   RBSr�
  G?Q�)$}�hMG?1�)$}�X   POSr�
  G?P�ƒ6BX   CCr�
  G?D�I��NG?!�)$}�X   ''r�
  G?:�=���X   WDTr�
  G?*�=���X   NNPSr�
  G?!�)$}�uj  j�
  �r�
  h h(h
c__builtin__
__main__
hNN}r�
  Ntr�
  Rr�
  �r�
  Rr�
  (X   VBDr�
  G?���Cm�X   VBNr�
  G?�sSކKX   POSr�
  G?�zE��h�G?����� �X   NNPr�
  G?�k����X   VBr�
  G?����bX   NNr�
  G?�8��^�X   RBr�
  G?���{u�GX   INr�
  G?��[:���X   MDr�
  G?V��{u�GX   CCr�
  G?|}��R��X   VBGr�
  G?����g�X   TOr�
  G?rGg��hMG?v��{u�GX   NNSr�
  G?w��+E&*X   oovr�
  G?Z�[:���X   DTr�
  G?�'M�8&X   JJr�
  G?�*�2�X   NNPSr�
  G?b�e�7Q�X   RBSr�
  G?^c���_X   JJSr�
  G?Nc���_X   CDr�
  G?�%	�ȟX   VBPr�
  G?^c���_X   ''r�
  G?>c���_X   JJRr�
  G?Nc���_X   WPr�
  G?>c���_X   VBZr�
  G?h���X   PRPr�
  G?R�e�7Q�NG?F��{u�GX   WDTr�
  G?>c���_X   WRBr�
  G?>c���_uj�
  j�  �r   h h(h
c__builtin__
__main__
hNN}r  Ntr  Rr  �r  Rr  (h�G?�iW�BX   WDTr  G?sp�Z�X   VBr  G?�k��y�[X   NNPr  G?��#�tFxX   DTr	  G?�A�pc$�X   PRP$r
  G?yE���QX   INr  G?�[�V�X   PRPr  G?cp�Z�X   VBGr  G?sp�Z�X   WPr  G?�	�P�X   RBr  G?�[�V�X   NNPSr  G?_��@�X   NNr  G?������X   JJr  G?�0(�X   CDr  G?_��@�X   NNSr  G?�S��p�X   JJRr  G?O��@�X   oovr  G?cp�Z�X   WRBr  G?gS��p�X   VBNr  G?WS��p�NG?O��@�X   CCr  G?O��@�X   ``r  G?WS��p�X   JJSr  G?O��@�uj�  h��r  h h(h
c__builtin__
__main__
hNN}r  Ntr  Rr  �r   Rr!  NG?�      sX   VBZr"  j�
  �r#  h h(h
c__builtin__
__main__
hNN}r$  Ntr%  Rr&  �r'  Rr(  (X   NNr)  G?�9�A̜�X   JJr*  G?�8��|�X   ``r+  G?v���i��X   JJSr,  G?���d���X   VBGr-  G?z���6��X   RBSr.  G?�k/���X   RBr/  G?u���X   NNPr0  G?·P��5X   NNSr1  G?�2�ФaX   oovr2  G?_�*��X   CDr3  G?s�
.�X   VBNr4  G?`h��5t�X   DTr5  G?Z��h ��X   JJRr6  G?f�ױS��X   PRPr7  G?"����<Sh�G?7p�9'�hX   WPr8  G?@h��5t�X   NNPSr9  G?U���X   VBPr:  G?,!	w�Z|X   VBr;  G?E���X   INr<  G?b����<SX   CCr=  G?2����<SX   TOr>  G?"����<SX   VBDr?  G?"����<SuX   WPr@  jF  �rA  h h(h
c__builtin__
__main__
hNN}rB  NtrC  RrD  �rE  RrF  (X   DTrG  G?�D"e���X   JJrH  G?��vh�L�X   NNPrI  G?�!.�f�X   CDrJ  G?��:ߖ)X   VBNrK  G?��Ki-��X   NNSrL  G?�&]���X   INrM  G?�'F���X   TOrN  G?_���X   PRPrO  G?��g1��sX   NNrP  G?��T�`X   VBGrQ  G?y#6�IX   VBDrR  G?Zu�,R�X   RBrS  G?�'F���X   RBSrT  G?�*�V�KX   PRP$rU  G?Zu�,R�X   VBrV  G?�*�V�KX   VBZrW  G?~m����hMG?E*�V�KX   ``rX  G?o���X   JJRrY  G?�.�f�D�X   JJSrZ  G?o���X   VBPr[  G?O���X   WPr\  G?O���X   NNPSr]  G?q2�vh�MX   oovr^  G?e*�V�KX   CCr_  G?O���X   RPr`  G?E*�V�KX   POSra  G?E*�V�KujF  jG  �rb  h h(h
c__builtin__
__main__
hNN}rc  Ntrd  Rre  �rf  Rrg  (X   VBGrh  G?z�<���X   NNri  G?�L.R��X   NNSrj  G?̌�~���X   CDrk  G?��V�q�X   VBZrl  G?gNKt�X   JJSrm  G?������X   JJrn  G?���&��?X   NNPro  G?�vl9�'gX   INrp  G?�XW����X   JJRrq  G?z�<���X   RBSrr  G?����O�X   RBrs  G?s�Y]<�X   ``rt  G?b��*QX   CCru  G?R��*QX   VBDrv  G?gNKt�X   NNPSrw  G?v#�wb@X   VBrx  G?`Pg�X   WPry  G?d���O�X   VBNrz  G?r��*QX   VBPr{  G?b��*QX   MDr|  G?R��*QX   oovr}  G?[��8�yX   DTr~  G?R��*QX   TOr  G?B��*Qh�G?B��*QX   POSr�  G?B��*QX   PRP$r�  G?B��*QujG  jh  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   NNSr�  G?��1��gX   NNr�  G?�������X   JJr�  G?������X   CCr�  G?�w�քX   INr�  G?�3O%���X   WPr�  G?qw�քX   CDr�  G?z3O%���X   DTr�  G?��1��gX   NNPr�  G?������X   TOr�  G?qw�քX   VBPr�  G?qw�քX   VBr�  G?�w�քX   VBNr�  G?z3O%���X   RPr�  G?z3O%���X   RBr�  G?z3O%���X   ``r�  G?�w�քX   POSr�  G?qw�քh�G?qw�քX   JJRr�  G?qw�քX   VBDr�  G?qw�քujh  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   INr�  G?�[E9�h�G?ԅ��B�hMG?�����X   TOr�  G?�(���X   VBPr�  G?�!d,��X   NNSr�  G?�����X   VBGr�  G?�|�.�q�X   VBNr�  G?�_���IvX   VBDr�  G?�����X   CCr�  G?��@�x5mX   NNr�  G?�#�[EX   VBZr�  G?�|�.�q�X   WDTr�  G?�*K��a�X   JJr�  G?�����X   ``r�  G?a����X   MDr�  G?��V�AX   RBSr�  G?a����X   RBr�  G?��j�(�X   oovr�  G?*K��a�X   ''r�  G?j��s��X   JJRr�  G?a����X   DTr�  G?*K��a�X   VBr�  G?�B�Y!dX   POSr�  G?j��s��X   WRBr�  G?a����X   WPr�  G?j��s��X   NNPr�  G?a����uj�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   PRPr�  G?�Y'�o�X   DTr�  G?��1S�<X   NNSr�  G?��.Y���X   JJr�  G?��/���X   INr�  G?��U�K�tX   NNPr�  G?�dgw� �X   WDTr�  G?������X   CDr�  G?�m(e�mX   VBGr�  G?�0�ƞ�X   NNr�  G?��D�SX   PRP$r�  G?�V���0X   JJSr�  G?S�����h�G?�b�|�oYX   WPr�  G?�/���X   RBr�  G?i5�첿�X   TOr�  G?W�Tm�C\X   WRBr�  G?l�ꍸ�X   JJRr�  G?pt��fvX   VBPr�  G?PΕ�!�2X   ``r�  G?b5"rQ�X   VBNr�  G?fh�����X   NNPSr�  G?L�ꍸ�X   oovr�  G?U;o�J~X   CCr�  G?6h�����NG?<�ꍸ�X   VBZr�  G?&h�����X   VBDr�  G?<�ꍸ�X   MDr�  G?&h�����uj�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (h�G?��uV��X   VBDr�  G?��@1L�X   INr�  G?��@��,*X   VBZr�  G?ɭQ��X   CDr�  G?`n��UX   VBr�  G?x�c��X   TOr�  G?����c^�X   RBr�  G?����D�hMG?x�c��X   MDr�  G?���$��X   VBPr�  G?�L�~T��X   WRBr�  G?h�c��X   VBGr�  G?|�L�~UX   NNr�  G?��L�~UX   CCr�  G?�|�U��X   JJRr�  G?`n��UX   DTr�  G?t���5�X   JJr�  G?����C��X   WPr�  G?`n��UX   NNSr�  G?h�c��X   oovr�  G?h�c��X   VBNr�  G?`n��UX   WDTr�  G?h�c��X   NNPr�  G?`n��UX   JJSr�  G?`n��UX   ``r�  G?t���5�uj�  h��r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (NG?��	Q��X   ``r�  G?�����+�X   ''r�  G?�����+�X   VBr   G?zP�XA�X   NNPr  G?q����+�uNh!�r  h h(h
c__builtin__
__main__
hNN}r  Ntr  Rr  �r  Rr  (X   NNr  G?�`��)	�X   POSr	  G?�R�ψ4X   VBZr
  G?��i��yX   VBDr  G?�}H��?�X   INr  G?���0i*�X   MDr  G?rJ0 �8X   NNPr  G?���MT�GX   RBr  G?��"4��hMG?�-�4��\h�G?E�&h�CX   CCr  G?�vm*�?X   NNSr  G?���)��IX   VBPr  G?u�$��@X   CDr  G?��Z"h]�X   WPr  G?th#56>X   JJr  G?�܁���X   oovr  G?�Yd1�oWX   VBGr  G?rJ0 �8X   WDTr  G?u�$��@X   DTr  G?���76Z�X   VBNr  G?RJ0 �8X   VBr  G?rJ0 �8X   WRBr  G?i�,�\NX   TOr  G?RJ0 �8X   NNPSr  G?`u��r2X   PRPr  G?th#56>X   PRP$r   G?RJ0 �8X   JJRr!  G?=C�36 ZX   ``r"  G?E�&h�CX   RBSr#  G?E�&h�CuX   PRP$r$  j3  �r%  h h(h
c__builtin__
__main__
hNN}r&  Ntr'  Rr(  �r)  Rr*  (X   INr+  G?��`v���X   NNr,  G?ݮ`v���X   NNPr-  G?��B�YX   JJSr.  G?��`v���X   NNSr/  G?�J3�)h�G?��`v���X   JJr0  G?�B�Y!dX   CCr1  G?��`v���X   VBGr2  G?��`v���hMG?��`v���uj3  j+  �r3  h h(h
c__builtin__
__main__
hNN}r4  Ntr5  Rr6  �r7  Rr8  (X   DTr9  G?�,�v�PX   NNPr:  G?�^~P��X   PRP$r;  G?��`�i��X   NNr<  G?��7�3�X   WRBr=  G?�6zt���X   PRPr>  G?�$(F޼X   WPr?  G?��ੳӥX   NNSr@  G?��[����X   CDrA  G?��ੳӥh�G?��ੳӥX   VBNrB  G?w$(F޼X   WDTrC  G?�$(F޼X   RBrD  G?sH�jdGX   JJrE  G?�h�!�e�X   INrF  G?����}Y1X   VBGrG  G?�։��X   ``rH  G?g$(F޼X   JJRrI  G?^�ੳӥX   TOrJ  G?^�ੳӥX   NNPSrK  G?^�ੳӥX   JJSrL  G?g$(F޼X   VBPrM  G?^�ੳӥX   VBDrN  G?^�ੳӥuj9  j  �rO  h h(h
c__builtin__
__main__
hNN}rP  NtrQ  RrR  �rS  RrT  (X   CDrU  G?b�N���KX   JJrV  G?��܆̐Bh�G?��"J~��X   NNSrW  G?�6�܆̐X   NNPrX  G?��N���KX   NNrY  G?�'R.�X   CCrZ  G?b�N���KX   RBr[  G?������6X   VBNr\  G?r�N���KX   TOr]  G?r�N���KX   INr^  G?��N���KX   WPr_  G?b�N���KX   VBr`  G?|`���9�X   NNPSra  G?b�N���KX   oovrb  G?b�N���Kuj  jU  �rc  h h(h
c__builtin__
__main__
hNN}rd  Ntre  Rrf  �rg  Rrh  (X   WPri  G?�      X   JJrj  G?�      ujU  ji  �rk  h h(h
c__builtin__
__main__
hNN}rl  Ntrm  Rrn  �ro  Rrp  (X   NNSrq  G?�z�G�{h�G?��Q��X   VBDrr  G?ۅ�Q�X   NNrs  G?�ffffffX   VBZrt  G?�z�G�{X   MDru  G?�z�G�{X   JJrv  G?�z�G�{X   NNPrw  G?�z�G�{X   RBrx  G?�z�G�{ujE  jV  �ry  h h(h
c__builtin__
__main__
hNN}rz  Ntr{  Rr|  �r}  Rr~  (X   NNr  G?��0�h)�X   JJr�  G?���}��;X   NNSr�  G?��e!���X   RBr�  G?a�����X   VBNr�  G?�?�]$ZX   INr�  G?�RO��mX   TOr�  G?��p��X   NNPr�  G?��p��X   VBDr�  G?a�����h�G?���7�X   VBGr�  G?~� ӢN�X   oovr�  G?q�����X   CCr�  G?�?�]$ZX   DTr�  G?a�����X   WPr�  G?jtI����X   CDr�  G?a�����X   ''r�  G?a�����hMG?jtI����X   NNPSr�  G?a�����X   VBr�  G?a�����X   VBPr�  G?a�����ujl  j
  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   INr�  G?�X   NNPr�  G?ˑ���X   CCr�  G?���X   POSr�  G?ũZ��Z�X   VBDr�  G?�YE�YE�h�G?�=��=��X   VBNr�  G?�����X   NNr�  G?�����X   RBr�  G?�X   NNSr�  G?�����X   TOr�  G?�PPX   VBr�  G?�����X   PRP$r�  G?o���� X   NNPSr�  G?uPPX   VBPr�  G?�a&a&X   MDr�  G?�a&a&hMG?��z�zX   JJr�  G?�����X   RBSr�  G?ePPX   VBZr�  G?�PPX   JJRr�  G?ePPX   PRPr�  G?ePPX   DTr�  G?zA�A�X   VBGr�  G?uPPNG?o���� X   ``r�  G?o���� X   oovr�  G?o���� X   CDr�  G?ePPuj.  j  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   NNPr�  G?���kC7�X   NNr�  G?�a@[�ݭX   JJr�  G?�s��JX   RBSr�  G?���kC7�X   NNSr�  G?�v�3|l�X   CDr�  G?���kC7�X   JJSr�  G?�)y�ri�X   NNPSr�  G?���kC7�X   VBGr�  G?���kC7�X   DTr�  G?���kC7�X   INr�  G?���kC7�uj�  jO  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   INr�  G?����_�\X   POSr�  G?��}+f�X   VBDr�  G?�(�o��X   NNr�  G?��g'�eh�G?�\v@(AjX   DTr�  G?�(�o��X   CCr�  G?����
X   NNPr�  G?ʻp��N�X   TOr�  G?������'X   NNSr�  G?�ީ��s�X   VBNr�  G?����*${X   WPr�  G?t �&^YQX   VBGr�  G?� �&^YQX   CDr�  G?�1����X   JJr�  G?�(�o��X   RBr�  G?�1����X   PRP$r�  G?~1����X   oovr�  G?�(�o��hMG?�(�o��X   MDr�  G?t �&^YQX   VBr�  G?�(�o��X   WDTr�  G?~1����X   PRPr�  G?~1����X   ``r�  G?t �&^YQX   VBPr�  G?t �&^YQX   NNPSr�  G?t �&^YQuX   JJr�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   NNr�  G?�%����X   JJr�  G?�Q�n��h�G?�G���X   INr�  G?���)�%X   CDr�  G?V�F���#X   VBDr�  G?t����X   NNSr�  G?�d@�F�X   VBNr�  G?�}�B��[X   NNPr�  G?��9A؆X   TOr�  G?�Ia/ú�X   WPr�  G?P{���>X   CCr�  G?�����X   VBGr�  G?l�ǥ�X   VBPr�  G?I�,?���X   JJSr�  G?CIa/ú�X   NNPSr�  G?v�F���#X   VBZr�  G?i�,?���X   PRP$r�  G?9�,?���X   RBr�  G?f�F���#hMG?a��k��wX   ''r�  G?p{���>X   VBr�  G?I�,?���X   DTr�  G?CIa/ú�NG?CIa/ú�X   WDTr�  G?CIa/ú�X   oovr�  G?CIa/ú�X   ``r�  G?CIa/ú�X   POSr�  G?CIa/ú�uX   VBr   h��r  h h(h
c__builtin__
__main__
hNN}r  Ntr  Rr  �r  Rr  (X   INr  G?Î8�8�h�G?�q�q�X   RPr  G?�����/hX   DTr	  G?�UUUUUUX   VBZr
  G?�B^З�&X   NNSr  G?|q�q�X   TOr  G?�q�q�X   VBNr  G?���%�	{X   VBDr  G?�%�	{B_X   ''r  G?r����/hX   VBr  G?�����/X   RBr  G?�З�%�	X   JJr  G?��q�rX   MDr  G?�����/X   JJRr  G?�����/hX   VBGr  G?��%�	{BhMG?r����/hX   VBPr  G?�UUUUUUX   oovr  G?�����/hX   JJSr  G?r����/hX   NNr  G?���%�	{X   WRBr  G?r����/hX   PRPr  G?|q�q�X   NNPr  G?r����/hX   WPr  G?|q�q�X   WDTr  G?r����/huh�j  �r  h h(h
c__builtin__
__main__
hNN}r   Ntr!  Rr"  �r#  Rr$  (X   DTr%  G?̳��?��X   NNr&  G?�E�t]FX   NNPr'  G?���|X   PRP$r(  G?�+qB�+X   JJr)  G?�שz��X   PRPr*  G?���0�X   VBGr+  G?��	O ��X   INr,  G?�+qB�+X   CDr-  G?���|X   WPr.  G?���0�X   NNSr/  G?�+qB�+h�G?�`1�`X   JJRr0  G?x��0�X   TOr1  G?���0�X   ``r2  G?��A)��X   VBNr3  G?��A)��X   VBDr4  G?���|X   RBr5  G?���0�hMG?��A)��X   WDTr6  G?x��0�uX   WDTr7  j+  �r8  h h(h
c__builtin__
__main__
hNN}r9  Ntr:  Rr;  �r<  Rr=  (X   VBDr>  G?�ffffffX   INr?  G?�������X   VBPr@  G?˻�����X   NNSrA  G?�X   VBNrB  G?�h�G?Ȉ�����X   MDrC  G?�333333X   VBZrD  G?�������X   PRP$rE  G?�X   NNrF  G?�UUUUUUX   oovrG  G?�X   VBGrH  G?�X   CCrI  G?�UUUUUUX   POSrJ  G?�X   DTrK  G?�������X   TOrL  G?�������X   VBrM  G?�X   RBrN  G?�������X   WDTrO  G?�uX   DTrP  j  �rQ  h h(h
c__builtin__
__main__
hNN}rR  NtrS  RrT  �rU  RrV  (X   JJSrW  G?�[b���+X   NNPrX  G?��I���X   JJrY  G?�&p�'�X   WPrZ  G?f���ُ	X   NNr[  G?�>B��IX   NNSr\  G?�v�!���X   VBNr]  G?r���5L�h�G?�.�bзX   INr^  G?�+(r%�X   RBSr_  G?x���JX   POSr`  G?����JhMG?�	n���X   VBDra  G?�i��}ъX   VBPrb  G?b���5L�X   WDTrc  G?^/��"X   CDrd  G?x���JX   CCre  G?��q�YX   NNPSrf  G?x���JX   TOrg  G?�	n���X   ``rh  G?V���ُ	X   VBZri  G?n/��"X   RBrj  G?^/��"X   VBGrk  G?f���ُ	X   DTrl  G?^/��"X   MDrm  G?N/��"X   oovrn  G?^/��"NG?N/��"X   ''ro  G?V���ُ	X   PRPrp  G?V���ُ	uj  jW  �rq  h h(h
c__builtin__
__main__
hNN}rr  Ntrs  Rrt  �ru  Rrv  (X   JJrw  G?��q�rX   NNSrx  G?ԟI��I�X   NNry  G?�������X   VBGrz  G?�X   RBr{  G?�X   INr|  G?�q�q�X   VBPr}  G?��l�lX   CDr~  G?��l�lujW  jw  �r  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   NNSr�  G?�A�j�p�X   NNr�  G?��k�QX   JJr�  G?���+(7X   NNPr�  G?�c��۵h�G?��L�x��X   VBNr�  G?oc��۵X   INr�  G?��v��X   VBGr�  G?w�L�x��X   TOr�  G?w�L�x��X   RBr�  G?���k�QhMG?oc��۵X   CCr�  G?oc��۵ujw  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   INr�  G?�����j�X   VBZr�  G?�<��X   VBDr�  G?��L;ˌ�h�G?�%��6�X   VBPr�  G?�0F�ZHX   VBNr�  G?�ռHVX   NNr�  G?�kϴ�p�hMG?�d#DpP�X   NNPr�  G?a.��@iX   TOr�  G?�Eq����X   MDr�  G?�$�gN�8X   RBr�  G?�Q��E�X   CCr�  G?�*�~BXX   ''r�  G?e�!����X   VBr�  G?����mQX   VBGr�  G?|�ׄ΋�X   JJr�  G?~5���X   POSr�  G?io��g�X   NNSr�  G?w �'�MX   WDTr�  G?��&��IX   DTr�  G?o�X��TNX   ``r�  G?F,>�D%X   WPr�  G?h�F��X   WRBr�  G?_
q�{�NG?F,>�D%X   JJSr�  G?:�=!�X   oovr�  G?a.��@iX   RPr�  G?F,>�D%X   RBSr�  G?F,>�D%X   JJRr�  G?L�ׄ΋�X   CDr�  G?1��eki�X   PRPr�  G?1��eki�X   NNPSr�  G?!��eki�X   PRP$r�  G?*�=!�ujP  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   NNPr�  G?�_��j��X   PRPr�  G?� 5���X   DTr�  G?�vL��X   VBNr�  G?��N���X   NNSr�  G?��3=��X   JJr�  G?�3s���X   WPr�  G?��Z��EX   TOr�  G?�{�4�JX   INr�  G?� 5���X   VBr�  G?w�Z��EX   NNr�  G?� 5���X   RBr�  G?��e9UX   NNPSr�  G?d))_";9X   ``r�  G?j�~�N�X   JJRr�  G?~=��X�X   CDr�  G?��~�N�X   oovr�  G?j�~�N�X   VBGr�  G?��Z��EX   RPr�  G?p���G1Zh�G?z�~�N�X   VBZr�  G?d))_";9X   RBSr�  G?d))_";9X   VBDr�  G?Z�~�N�X   JJSr�  G?d))_";9X   POSr�  G?Z�~�N�uj�  j�
  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   INr�  G?����}�^h�G?�τ���LX   VBDr�  G?\�����X   TOr�  G?�m�&кX   DTr�  G?������X   NNSr�  G?z���N�X   VBNr�  G?�τ���LX   RBr�  G?��g�pX   VBGr�  G?���[��X   JJr�  G?sU5P�X   NNr�  G?�*J���X   ``r�  G?SU5P�X   RPr�  G?p�g�pX   PRPr�  G?\�����X   CDr�  G?cU5P�X   VBr�  G?SU5P�X   NNPr�  G?p�g�pNG?cU5P�X   WRBr�  G?SU5P�hMG?SU5P�X   VBZr�  G?SU5P�X   CCr�  G?SU5P�uj�
  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   PRP$r�  G?�G���X   WPr�  G?�"�7t�"h�G?��|t0X   DTr�  G?�b�xX   WDTr�  G?��C�2�+X   NNPr�  G?ƫ��Q��X   CDr�  G?��vJ(X   NNr�  G?�����-�X   VBGr�  G?���|tX   PRPr�  G?xӁ����X   INr�  G?���ͳ�X   NNSr�  G?�_o��BX   JJr�  G?�{���X   WRBr�  G?t�	�+�OX   ``r�  G?g�㠐q~X   VBDr�  G?N�1�X   NNPSr   G?I��Ӂ�X   TOr  G?i&�gђX   RBr  G?v?1�9dX   VBNr  G?Y��Ӂ�X   JJRr  G?b�C�2�+X   JJSr  G?g�㠐q~hMG?T��vJX   CCr  G?U짨Ma_X   VBr  G?$��vJX   oovr  G?P����X   VBZr	  G?I��Ӂ�X   ''r
  G?$��vJX   VBPr  G?4��vJNG?B/��A!X   MDr  G?$��vJuj�  j,  �r  h h(h
c__builtin__
__main__
hNN}r  Ntr  Rr  �r  Rr  (X   NNr  G?��k�egX   POSr  G?}������X   VBDr  G?�ھ�P^h�G?�ziae��X   INr  G?�V8jq�dX   TOr  G?�m$�6�X   CDr  G?a���X   RBr  G?������X   JJr  G?�(�5�2�X   VBNr  G?��:14hMG?�{y�!�X   NNSr  G?�8jq�c�X   WDTr  G?���A��X   CCr  G?�j�%Av�X   DTr  G?��;��X   WRBr   G?uI���T�X   JJRr!  G?Y�����X   NNPr"  G?�{y�!��X   VBZr#  G?����X   VBGr$  G?��A��X   VBr%  G?wj�%Av�NG?s(�5�2�X   PRP$r&  G?eI���T�X   WPr'  G?}������X   oovr(  G?a���X   ''r)  G?a���X   MDr*  G?m������X   PRPr+  G?uI���T�X   VBPr,  G?a���X   ``r-  G?Q���uX   INr.  jJ  �r/  h h(h
c__builtin__
__main__
hNN}r0  Ntr1  Rr2  �r3  Rr4  (X   NNPr5  G?�U��E�h�G?���	�xX   NNr6  G?��%���}X   CDr7  G?��|�SX   INr8  G?���G�!X   NNSr9  G?�`iˣm�X   ``r:  G?l����MX   PRP$r;  G?��k�U�X   DTr<  G?���'�X   JJr=  G?����k�X   VBNr>  G?���'�X   TOr?  G?�1�T�v	X   RPr@  G?���[��X   WPrA  G?�p�,�yX   WRBrB  G?{)�;T�X   POSrC  G?Q'��"�X   WDTrD  G?i��{���X   CCrE  G?�r��t?�X   PRPrF  G?���'�hMG?os�z��X   MDrG  G?os�z��X   VBPrH  G?t�|�SX   VBGrI  G?r���:�X   RBrJ  G?�p�,�yX   ''rK  G?V����qX   JJRrL  G?r���:�X   VBDrM  G?v����qX   oovrN  G?i��{���X   VBrO  G?d�|�SX   VBZrP  G?\����MX   NNPSrQ  G?F����quX   VBDrR  h��rS  h h(h
c__builtin__
__main__
hNN}rT  NtrU  RrV  �rW  RrX  (NG?�����X�X   ''rY  G?T��Q��.X   INrZ  G?K]¥@>uj	  jN  �r[  h h(h
c__builtin__
__main__
hNN}r\  Ntr]  Rr^  �r_  Rr`  (X   NNra  G?�UUUUUUX   VBNrb  G?�a�a�X   NNSrc  G?�I$�I$�X   JJrd  G?�a�a�ujN  ja  �re  h h(h
c__builtin__
__main__
hNN}rf  Ntrg  Rrh  �ri  Rrj  (X   RBrk  G?�X   INrl  G?ӳ�����h�G?�������X   POSrm  G?�X   TOrn  G?�X   NNSro  G?�������X   CCrp  G?�X   WRBrq  G?pX   NNrr  G?�������X   VBDrs  G?�X   MDrt  G?�X   VBZru  G?�X   VBNrv  G?�X   VBGrw  G?�hMG?�X   NNPrx  G?�X   VBPry  G?�X   VBrz  G?xX   ''r{  G?pX   JJr|  G?�X   WPr}  G?xX   PRPr~  G?pX   PRP$r  G?puja  jk  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   VBDr�  G?ŕ<
��X   VBZr�  G?��v�&��X   INr�  G?��\��X   WPr�  G?\�Ak=<�X   RBr�  G?�.����hMG?|�Ak=<�h�G?����X   TOr�  G?�����0�X   VBNr�  G?�Xk��R&X   VBPr�  G?��$%
t�X   VBGr�  G?��Ak=<�X   VBr�  G?���m�{X   oovr�  G?|�Ak=<�X   NNr�  G?��H�E�X   JJr�  G?��=ՕX   DTr�  G?�׬\X   WRBr�  G?zI{����X   NNSr�  G?�׬\X   ''r�  G?S+��}�X   MDr�  G?g嶄]3X   NNPr�  G?l�Ak=<�X   CCr�  G?zI{����X   PRPr�  G?\�Ak=<�X   CDr�  G?c+��}�NG?c+��}�X   JJRr�  G?\�Ak=<�X   JJSr�  G?\�Ak=<�X   ``r�  G?S+��}�ujk  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   INr�  G?�:��ˑX   NNPr�  G?���e�]�X   DTr�  G?ӄ̒:�X   PRPr�  G?�S` �X   WDTr�  G?[�\f�h�X   VBNr�  G?��$�F�X   WPr�  G?�[�����X   TOr�  G?�z��^CX   NNSr�  G?��� $�{X   PRP$r�  G?}�$�F�h�G?�8p+��X   JJr�  G?�u�VX   NNr�  G?�3�9���X   RPr�  G?�V=���cX   RBr�  G?�[�����X   JJSr�  G?f�� $�{X   WRBr�  G?t�L��oX   VBGr�  G?t�L��oX   ``r�  G?k�\f�h�X   JJRr�  G?[�\f�h�X   CCr�  G?v�� $�{X   CDr�  G?y6��[��hMG?k�\f�h�X   ''r�  G?bV=���cX   VBr�  G?f�� $�{X   oovr�  G?bV=���cX   NNPSr�  G?[�\f�h�uj�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   WPr�  G?�      X   DTr�  G?�      X   VBGr�  G?�      X   NNSr�  G?�      h�G?�      X   NNPr�  G?�      X   CDr�  G?�      uj-	  h��r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (NG?��fffffX   WPr�  G?9������X   ''r�  G?9������X   NNr�  G?9������uNh"�r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   POSr�  G?����ȫ)X   NNr�  G?�!�����X   VBDr�  G?���X��X   CCr�  G?������X   INr�  G?�!�����X   VBZr�  G?���%��X   VBNr�  G?}�����X   NNSr�  G?�ÁK�X   NNPr�  G?������X   MDr�  G?�.zw��X   DTr�  G?ʾWm0X   CDr�  G?��5?rZX   VBGr�  G?���- �hMG?��_�dVX   RBr�  G?q���ȫ)X   TOr�  G?������X   WDTr�  G?���k�9�NG?q���ȫ)X   PRP$r�  G?g��k�9�X   WRBr�  G?g��k�9�uh"j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   NNr�  G?�<g��4X   JJr�  G?��<g��X   CDr�  G?�B(E�X   JJSr�  G?�      X   NNSr�  G?��p.�X   NNPr�  G?�Øsa�X   RBSr�  G?�SjmM��h�G?�.��X   VBDr�  G?�B(E�X   POSr�  G?qB(E�X   WPr�  G?g�\�pX   INr�  G?|Øsa�X   VBZr�  G?W�\�pX   WRBr�  G?W�\�pX   ``r�  G?lØsa�X   RBr�  G?g�\�pX   VBNr   G?y�<g��X   VBGr  G?g�\�pX   VBPr  G?qB(E�hMG?g�\�pX   oovr  G?aB(E�X   JJRr  G?W�\�pX   MDr  G?W�\�pX   TOr  G?aB(E�X   DTr  G?qB(E�X   VBr  G?g�\�pX   CCr	  G?qB(E�X   ''r
  G?aB(E�uX   DTr  j  �r  h h(h
c__builtin__
__main__
hNN}r  Ntr  Rr  �r  Rr  (X   NNr  G?��쳍FDX   VBGr  G?�m�D<��X   DTr  G?|%��J�h�G?�I[)yޅX   VBPr  G?��]�'W�X   VBNr  G?����@ӊX   INr  G?�:�iW�X   NNPr  G?���BX   WDTr  G?�ky��dX   VBDr  G?�N����X   MDr  G?w�%QZOhMG?�t���i!X   NNSr  G?�����NX   TOr  G?��v��X   CCr  G?�Ȏr�%X   PRPr  G?tx�E�>X   VBr   G?w�%QZOX   RBr!  G?�ب	a�`X   WPr"  G?�|m���ZX   JJSr#  G?b����NX   POSr$  G?�t���i!X   JJr%  G?�Ȏr�%X   WRBr&  G?kK�\�~�X   oovr'  G?W�%QZOX   VBZr(  G?w�%QZOX   RPr)  G?Q?:�^X   JJRr*  G?;K�\�~�X   ``r+  G?i���)�X   CDr,  G?W�%QZOX   ''r-  G?[K�\�~�NG?Q?:�^X   RBSr.  G?;K�\�~�X   PRP$r/  G?;K�\�~�uj  j  �r0  h h(h
c__builtin__
__main__
hNN}r1  Ntr2  Rr3  �r4  Rr5  (X   INr6  G?�*�r���h�G?��M"�X   VBDr7  G?���dC�
X   NNSr8  G?�Ռ�"`\X   TOr9  G?�z��u19X   NNr:  G?��:U��-X   VBZr;  G?�:�G�PX   VBNr<  G?� K �X   VBr=  G?y B�\s�X   JJr>  G?����}DX   VBPr?  G?���9���X   DTr@  G?��2 �V�X   ''rA  G?tՌ�"`\X   CCrB  G?�
�*�sX   RBrC  G?����MX   VBGrD  G?}*�r���X   PRPrE  G?tՌ�"`\X   NNPrF  G?� B�\s�X   CDrG  G?`���MX   MDrH  G?}*�r���X   WDTrI  G?p���MhMG?}*�r���NG?p���MX   WPrJ  G?`���MX   WRBrK  G?p���MX   ``rL  G?`���MX   POSrM  G?`���MuX   WPrN  j  �rO  h h(h
c__builtin__
__main__
hNN}rP  NtrQ  RrR  �rS  RrT  (X   NNrU  G?�����/hh�G?�����/hX   JJrV  G?Ǵ%�	{BX   NNPrW  G?�����/hX   INrX  G?�����/huX   NNPrY  jm  �rZ  h h(h
c__builtin__
__main__
hNN}r[  Ntr\  Rr]  �r^  Rr_  (X   VBDr`  G?�+�:i�.X   INra  G?��-CͪX   VBPrb  G?���Xv�X   VBZrc  G?��y�TT�X   VBrd  G?�W& �LAX   NNSre  G?b�s��X   oovrf  G?r�s��X   RBrg  G?���Pc+cX   TOrh  G?�G�N�nX   JJri  G?�(a����X   VBNrj  G?��ؾ�}h�G?�짉LHX   NNrk  G?�i^+�X   CDrl  G?h
��a{X   VBGrm  G?��7�R�(X   DTrn  G?���Pc+cX   WRBro  G?b�s��X   NNPrp  G?n%��9�X   NNPSrq  G?X
��a{X   JJRrr  G?h
��a{NG?X
��a{X   MDrs  G?X
��a{hMG?b�s��X   CCrt  G?n%��9�X   JJSru  G?X
��a{uX   NNPrv  j
  �rw  h h(h
c__builtin__
__main__
hNN}rx  Ntry  Rrz  �r{  Rr|  (X   DTr}  G?���|#�X   NNPr~  G?�>��L�X   RBr  G?�6���|`X   PRP$r�  G?�4&}5WX   JJSr�  G?s�*�`X   VBNr�  G?�}���ɶX   NNr�  G?��\/
�jh�G?���@&�X   INr�  G?�H�4cO�X   WPr�  G?�KP�)u}X   VBr�  G?���9��X   JJr�  G?�d���sX   oovr�  G?x��7�i}X   PRPr�  G?�~(���X   NNSr�  G?��\/
�jX   WRBr�  G?���7�i}X   RPr�  G?s�*�`X   WDTr�  G?�'�$Y��X   ``r�  G?q4&}5WX   TOr�  G?�ۦ1.5�X   VBDr�  G?��*�`X   VBGr�  G?��\/
�jhMG?j�;�6�X   JJRr�  G?|��@&�X   CDr�  G?���3Q�sX   POSr�  G?Ni@DlКX   VBPr�  G?x��7�i}X   CCr�  G?V��3Q�sX   VBZr�  G?v��3Q�sX   RBSr�  G?^i@DlКX   MDr�  G?V��3Q�suX   NNr�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   WRBr�  G?v�:��zX   INr�  G?�»!���h�G?�I$�I$�X   TOr�  G?����l�X   JJr�  G?���/9X   NNr�  G?�� Ŕ�X   NNSr�  G?���@e�X   CCr�  G?�,+��X   VBGr�  G?z��`jc�X   NNPr�  G?���"���hMG?r��ip�cX   VBPr�  G?ne���MkX   VBZr�  G?���/9X   VBDr�  G?�,+��X   PRPr�  G?f�:��zX   RBr�  G?�I�(ؔX   RPr�  G?f�:��zX   ``r�  G?��:��zX   VBr�  G?r��ip�cX   VBNr�  G?���ip�cX   CDr�  G?^e���MkNG?f�:��zX   WDTr�  G?f�:��zX   ''r�  G?^e���MkX   NNPSr�  G?^e���Mkuj�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   NNPr�  G?�������X   PRPr�  G?�������X   VBDr�  G?�333333X   TOr�  G?�������X   JJr�  G?�������h�G?�333333X   INr�  G?�������X   WPr�  G?�������X   DTr�  G?�������X   NNr�  G?�������X   NNSr�  G?�������X   RBr�  G?�������X   VBGr�  G?�ffffffX   VBNr�  G?�������X   VBZr�  G?�������uj�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   VBDr�  G?��CV��X   NNPr�  G?�41�o�<X   VBZr�  G?��,��X   NNr�  G?�ڷ��CX   VBPr�  G?��CV��X   PRPr�  G?��,��X   CCr�  G?�ڷ��CX   POSr�  G?�'�Yy�RX   NNSr�  G?��CV��X   MDr�  G?��,��X   VBr�  G?��,��X   CDr�  G?��CV��X   RBr�  G?��,��hMG?��CV��uj�  j,  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   NNr�  G?�h1���X   INr�  G?����%B�X   JJr�  G?����%B�X   NNSr�  G?�73��|4X   NNPr�  G?���Ĩ]�h�G?v�h1��X   NNPSr�  G?����%B�X   VBZr�  G?v�h1��X   PRPr�  G?v�h1��X   VBDr�  G?��h1��hMG?v�h1��X   RBr�  G?��h1��X   CDr�  G?����%B�X   DTr�  G?v�h1��X   TOr�  G?v�h1��X   VBGr�  G?v�h1��uj  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   INr�  G?��.���X   WPr�  G?���Fl�X   WRBr�  G?���Fl�h�G?�`��a�X   TOr�  G?���|�/X   VBGr�  G?}$9y8v/X   NNPr�  G?���,�tX   DTr�  G?��a���X   RPr�  G?��ַY>�X   RBr   G?�?�=�+�X   NNr  G?�0��^X   PRPr  G?]$9y8v/X   JJRr  G?P0��^X   VBNr  G?�T����X   JJr  G?�3��qS�hMG?~®q��2X   PRP$r  G?V�e�+�%X   NNSr  G?p��1`�X   VBDr  G?]$9y8v/X   CDr	  G?Y�O�20*X   JJSr
  G?Sm{�%� X   CCr  G?u�+�X�X   ``r  G?]$9y8v/X   oovr  G?Y�O�20*X   MDr  G?P0��^NG?Sm{�%� X   WDTr  G?Cm{�%� X   ''r  G?V�e�+�%X   POSr  G?Cm{�%� X   VBZr  G?9�O�20*X   VBPr  G?9�O�20*uX   VBr  h��r  h h(h
c__builtin__
__main__
hNN}r  Ntr  Rr  �r  Rr  (X   NNr  G?�F�`FX   VBr  G?�B9$#�Bh�G?�Z���[X   DTr  G?���� X   NNPr  G?�11�X   RBr  G?���
h�X   VBGr   G?���
h�X   NNSr!  G?�*"�*X   JJr"  G?�*"�*X   INr#  G?���_,�X   ``r$  G?X8��8X   WPr%  G?�vAwdvX   PRP$r&  G?���
h�X   NNPSr'  G?X8��8X   CDr(  G?r*"�*X   TOr)  G?b*"�*X   PRPr*  G?�*"�*X   WRBr+  G?u1S1X   WDTr,  G?X8��8X   CCr-  G?X8��8X   JJRr.  G?X8��8X   oovr/  G?X8��8uh�j  �r0  h h(h
c__builtin__
__main__
hNN}r1  Ntr2  Rr3  �r4  Rr5  (X   INr6  G?�U�)�k�X   NNSr7  G?�N���Oh�G?�y�y�X   NNPr8  G?��8�8X   CCr9  G?�N���OX   DTr:  G?�t�{���X   NNr;  G?��Z�w�LX   VBNr<  G?�t�{���hMG?�n3��JX   PRPr=  G?wg��4��X   VBZr>  G?�N���OX   WPr?  G?wg��4��X   JJr@  G?��8�8X   ''rA  G?o5&����X   VBGrB  G?�g��4��X   RBrC  G?5&����X   MDrD  G?o5&����X   POSrE  G?��8�8X   VBDrF  G?o5&����X   PRP$rG  G?5&����X   VBrH  G?5&����X   TOrI  G?5&����X   WDTrJ  G?o5&����X   RPrK  G?o5&����X   CDrL  G?wg��4��X   ``rM  G?o5&����uX   POSrN  jO  �rO  h h(h
c__builtin__
__main__
hNN}rP  NtrQ  RrR  �rS  RrT  (X   NNrU  G?��.��X   NNSrV  G?�E�t]FX   WPrW  G?�E�t]FX   NNPrX  G?�t]E�tX   INrY  G?�E�t]FX   VBNrZ  G?�E�t]FX   WRBr[  G?�E�t]FX   RPr\  G?�E�t]FuX   TOr]  j  �r^  h h(h
c__builtin__
__main__
hNN}r_  Ntr`  Rra  �rb  Rrc  (X   NNrd  G?����l�X   JJre  G?��1&�yX   NNSrf  G?�z�G�{X   DTrg  G?��1&�yX   NNPrh  G?�z�G�{X   VBri  G?��t�j~�X   CDrj  G?�bM���X   RBrk  G?��t�j~�X   INrl  G?�bM���uj�  j�  �rm  h h(h
c__builtin__
__main__
hNN}rn  Ntro  Rrp  �rq  Rrr  (X   JJrs  G?�i:E�X   NNrt  G?�j�+���hMG?�i:E�X   NNSru  G?� �I��)h�G?�j�+���X   TOrv  G?��P �JX   INrw  G?�=@d��'X   NNPrx  G?�ؼw\��X   DTry  G?�ؼw\��X   MDrz  G?� �I��)X   CCr{  G?�������NG?� �I��)X   VBr|  G?� �I��)X   NNPSr}  G?� �I��)uj/  j�  �r~  h h(h
c__builtin__
__main__
hNN}r  Ntr�  Rr�  �r�  Rr�  (X   VBDr�  G?�',��[h�G?�N�,V?X   TOr�  G?�� M��`X   INr�  G?� M��_�hMG?�8{�}��X   VBPr�  G?�KO����X   WPr�  G?m',��[X   VBr�  G?��>@���X   RBr�  G?��jI}k3X   VBNr�  G?��G|ϷX   NNr�  G?��az�DTX   VBGr�  G?�KO����X   CCr�  G?�',��[X   DTr�  G?xKO����X   RPr�  G?xKO����X   oovr�  G?}',��[X   JJr�  G?������X   POSr�  G?sos��X   MDr�  G?�os��X   VBZr�  G?xKO����X   NNSr�  G?xKO����X   NNPr�  G?m',��[NG?m',��[X   WRBr�  G?xKO����X   JJRr�  G?cos��X   CDr�  G?cos��X   PRPr�  G?cos��X   ``r�  G?sos��uNh#�r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   WDTr�  G?�      X   VBDr�  G?�      X   VBPr�  G?�      X   VBZr�  G?�      X   MDr�  G?�      X   WPr�  G?�      uh#j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   NNr�  G?�t]E�tX   VBDr�  G?�t]E�tX   VBZr�  G?�t]E�tX   VBPr�  G?�E�t]FuX   NNPr�  h|�r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   NNr�  G?ڦ�N&�X   CDr�  G?��Y[fX   NNPr�  G?��\�*��X   JJSr�  G?�=2��vX   RBr�  G?��CΔԝX   RBSr�  G?�=2��vX   JJr�  G?˹��� xX   VBGr�  G?rcir�X   INr�  G?��CΔԝX   NNSr�  G?��CΔ�X   ``r�  G?��CΔ�X   VBPr�  G?��CΔԝX   VBr�  G?k�+�#X   VBDr�  G?k�+�#X   VBNr�  G?��CΔ�X   WPr�  G?bcir�X   DTr�  G?k�+�#X   VBZr�  G?bcir�X   NNPSr�  G?v�CΔԝX   oovr�  G?bcir�uNh$�r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   NNr�  G?����X   CDr�  G?�!m9M3X   JJr�  G?�rV{�o�X   NNPr�  G?���@��oX   VBPr�  G?�H�&3wX   INr�  G?���xp{X   VBZr�  G?�mL#��X   VBDr�  G?�3����X   RBr�  G?���xp{X   MDr�  G?u9	H��X   NNSr�  G?�)bk���X   CCr�  G?iw���X   PRPr�  G?`�m��s"X   JJSr�  G?`�m��s"X   DTr�  G?`�m��s"X   WDTr�  G?`�m��s"uX   NNr�  j�	  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (h�G?҄��֚�X   NNr�  G?Ǳ��T�X   VBZr�  G?���Zj��X   NNSr�  G?���Zj��X   INr�  G?�T�_�#�X   TOr�  G?�%	��5X   JJr�  G?�;�6w�mhMG?����֚�X   CCr�  G?���p4JX   NNPr�  G?������ X   VBDr�  G?���p4JX   ''r�  G?qn�BsyX   WRBr�  G?qn�BsyX   RBr�  G?�n�BsyX   VBr�  G?qn�BsyX   POSr�  G?�n�BsyX   VBNr�  G?�Ɉ+�WNG?�n�BsyX   MDr�  G?�Ɉ+�WX   WDTr�  G?qn�BsyX   JJRr�  G?�Ɉ+�WX   WPr�  G?qn�BsyX   CDr�  G?qn�BsyuX   NNPr�  h~�r   h h(h
c__builtin__
__main__
hNN}r  Ntr  Rr  �r  Rr  (X   PRPr  G?�W����MX   RBr  G?�:�[W��X   PRP$r  G?�:�[W��X   DTr	  G?�6�@�X   VBDr
  G?�	�r-��X   CDr  G?��V��X   INr  G?�:�[W��X   NNPr  G?�ι�h�G?�	�r-��X   JJr  G?�m^�ǃX   VBGr  G?�Ӈ���X   VBZr  G?�:�[W��X   NNr  G?��V��X   TOr  G?��V��X   VBNr  G?�:�[W��X   NNSr  G?��V��X   MDr  G?�:�[W��X   VBr  G?�:�[W��uX   INr  j�  �r  h h(h
c__builtin__
__main__
hNN}r  Ntr  Rr  �r  Rr  (X   CDr  G?��� �<X   DTr  G?�sF\їX   ``r   G?m�|A�X   NNPr!  G?�����!X   INr"  G?�7dM�vX   PRP$r#  G?�5�yC^X   NNr$  G?�Jڒ���X   NNSr%  G?��tŝ1X   VBGr&  G?�ї4e�h�G?�vDݑ7X   WRBr'  G?t��=aOXX   PRPr(  G?���X   JJSr)  G?w��@X   JJr*  G?�w��X   WPr+  G?�5�yC^X   CCr,  G?pw��|X   oovr-  G?g��@X   WDTr.  G?pw��|X   VBZr/  G?G��@X   JJRr0  G?W��@X   NNPSr1  G?G��@X   RBr2  G?d��=aOXX   TOr3  G?j򆼡�(X   VBNr4  G?Q�}�phMG?G��@uj  j�
  �r5  h h(h
c__builtin__
__main__
hNN}r6  Ntr7  Rr8  �r9  Rr:  (h�G?̾�oh �X   VBDr;  G?�eJ%��X   INr<  G?��:[�X   WRBr=  G?}�E���X   TOr>  G?�?:��X   VBZr?  G?��1�2X   MDr@  G?����eX   PRPrA  G?W��]d�X   NNPrB  G?�g��ۺX   WPrC  G?��_�|�X   VBNrD  G?���ː��X   WDTrE  G?���]d�X   VBPrF  G?�T�\	`[hMG?�.cpd�;X   RBrG  G?��f�/!X   VBGrH  G?��1�2X   NNSrI  G?y�dMz��X   DTrJ  G?��_�|�X   VBrK  G?}�E���X   ''rL  G?_�g��ۺX   NNrM  G?����eX   JJrN  G?���]d�X   CCrO  G?���U@GX   JJRrP  G?c�`�#)UX   oovrQ  G?g��]d�X   POSrR  G?c�`�#)UNG?W��]d�X   RBSrS  G?O�g��ۺX   CDrT  G?W��]d�X   ``rU  G?W��]d�uj�
  h��rV  h h(h
c__builtin__
__main__
hNN}rW  NtrX  RrY  �rZ  Rr[  (NG?��x�ۄIh�G?MBS^�X   WPr\  G?'he�K@�X   ''r]  G?Q�Le8pxX   ``r^  G?D{Y �،X   WRBr_  G?'he�K@�X   DTr`  G?'he�K@�X   NNPra  G?'he�K@�X   NNSrb  G?'he�K@�ujK  hM�rc  h h(h
c__builtin__
__main__
hNN}rd  Ntre  Rrf  �rg  Rrh  (X   WPri  G?�ۀ�69ZX   CDrj  G?��_i�UX   NNPrk  G?���/��hX   WRBrl  G?��`t�LX   WDTrm  G?�kg�oX   VBGrn  G?���@�X   VBNro  G?}2��>X   DTrp  G?�vZ����X   INrq  G?��"iQہX   VBDrr  G?�Hx���X   RBrs  G?}2��>X   NNSrt  G?��/r.�X   TOru  G?i�+FcX   NNrv  G?���N���X   JJrw  G?��`t�LX   oovrx  G?i�+FcX   CCry  G?���Eݖ�X   VBZrz  G?t��N���X   PRPr{  G?i�+FcX   VBPr|  G?p�/r.�X   RBSr}  G?`�/r.�hMG?`�/r.�X   NNPSr~  G?`�/r.�X   JJRr  G?`�/r.�uj�  j  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   NNr�  G?���\���X   DTr�  G?��"N&*X   NNPr�  G?�Kx~폧X   NNSr�  G?�p���C�X   INr�  G?�M/�ގX   TOr�  G?�rKx~�X   WRBr�  G?{q���k4h�G?�q���k4X   JJr�  G?���(��X   WPr�  G?�n4P��X   RBr�  G?�n4P��X   PRPr�  G?�q���k4X   RPr�  G?��9��gX   VBNr�  G?�LT�X   VBGr�  G?�q���k4X   PRP$r�  G?���Ռ8�X   JJRr�  G?kq���k4X   VBr�  G?t�9��gX   CDr�  G?�'� X   CCr�  G?��9��gX   VBDr�  G?{q���k4X   WDTr�  G?�'� X   VBZr�  G?t�9��gX   VBPr�  G?kq���k4uX   NNSr�  j  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   NNr�  G?�m�@�h�G?|X��I�X   NNSr�  G?�͂6�UX   JJr�  G?�%4CRapX   INr�  G?�X��I�X   NNPr�  G?�͂6�UX   VBDr�  G?�X��I�X   VBGr�  G?�Bo���$X   VBNr�  G?�X��I�X   VBPr�  G?��k.�X   RBSr�  G?�X��I�X   NNPSr�  G?|X��I�X   RBr�  G?|X��I�X   JJSr�  G?|X��I�X   VBZr�  G?|X��I�uX   NNPr�  h�r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   NNPr�  G?��O�jxX   WDTr�  G?u"��=�fX   VBr�  G?�`*E7�{X   VBGr�  G?u"��=�fX   NNr�  G?�����U�X   WPr�  G?�1#�g�h�G?��}�pX   PRP$r�  G?��|���X   DTr�  G?�'��B�kX   CDr�  G?p�|���X   WRBr�  G?u"��=�fX   NNSr�  G?i\��w�X   CCr�  G?`�|���X   RBr�  G?}��8�`�X   INr�  G?y\��w�X   PRPr�  G?i\��w�X   JJr�  G?}��8�`�X   NNPSr�  G?`�|���uhj�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   CCr�  G?���!�@X   POSr�  G?���(&�X   RBr�  G?w0�rh�G?Ճa�u�2X   INr�  G?�4aF�wKX   NNPr�  G?�k�S��TX   VBr�  G?t���N#fX   TOr�  G?��q��O�hMG?����|ytX   WPr�  G?rkY�~X[X   VBDr�  G?�kY�~X[X   WRBr�  G?bkY�~X[X   VBNr�  G?��zu��X   NNr�  G?������X   NNSr�  G?�%j0�X   NNPSr�  G?k�y���X   VBGr�  G?�zP�U�X   PRPr�  G?bkY�~X[X   VBZr�  G?rkY�~X[X   ''r�  G?[�y���X   DTr�  G?k�y���X   JJr�  G?}�q��O�X   CDr�  G?�0�rX   WDTr�  G?g0�rX   oovr�  G?bkY�~X[NG?p�q��PX   MDr�  G?bkY�~X[X   ``r�  G?[�y���X   VBPr�  G?RkY�~X[X   JJRr�  G?RkY�~X[uj�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   VBr�  G?��\�pX   INr�  G?�"�P�BX   VBDr�  G?��$o8��X   DTr�  G?�L�A2�X   NNr�  G?�-L�A3X   TOr�  G?��\�phMG?���z��X   PRPr�  G?���z��h�G?�ذkb��X   RBr�  G?�lX5�aX   NNSr�  G?��\�pX   VBGr�  G?���z��X   JJr�  G?��v�1�X   VBNr�  G?��nC�X   VBZr�  G?��\�pX   MDr�  G?��\�pX   oovr�  G?~��z��X   NNPr   G?�ذkb��X   CDr  G?~��z��X   VBPr  G?���z��X   WPr  G?�-L�A3X   JJRr  G?~��z��uj�  j�  �r  h h(h
c__builtin__
__main__
hNN}r  Ntr  Rr  �r	  Rr
  (X   PRPr  G?�v[R��h�G?��5���X   WDTr  G?j_�,�KX   JJr  G?�b���BDX   DTr  G?�sc��*X   INr  G?�$�J�X   NNr  G?��\OȜ�X   PRP$r  G?�_�,�KX   VBNr  G?�Q�5>y�X   NNPr  G?�����݌X   TOr  G?�L(8���X   WPr  G?�$�J�X   NNSr  G?�e��F9	X   RPr  G?���!���X   RBr  G?��';�X   JJRr  G?w����݌X   VBDr  G?e��o�X   VBGr  G?w����݌X   VBr  G?z_�,�KhMG?u��o�X   WRBr  G?�$�J�X   CDr  G?j_�,�KX   CCr  G?z_�,�KX   oovr   G?e��o�X   ``r!  G?o�Si'fX   MDr"  G?U��o�X   ''r#  G?_�Si'fX   NNPSr$  G?U��o�uX   NNPr%  jo  �r&  h h(h
c__builtin__
__main__
hNN}r'  Ntr(  Rr)  �r*  Rr+  (hMG?�ҶI�h�G?�S�K�X   NNr,  G?���/�T�X   CCr-  G?�Qz��;OX   NNPSr.  G?XA/.��X   NNPr/  G?���j~3X   INr0  G?��\H�X   WRBr1  G?u9	H��X   VBDr2  G?��s���X   NNSr3  G?�v��}��NG?xA/.��X   ``r4  G?hA/.��X   MDr5  G?b0�cV�X   JJr6  G?�IU��.X   VBZr7  G?���p-z8X   VBNr8  G?���V3ZX   VBGr9  G?xA/.��X   POSr:  G?u9	H��X   RBr;  G?���p-z8X   CDr<  G?�Qz��;OX   TOr=  G?��;��|X   VBPr>  G?xA/.��X   oovr?  G?�A/.��X   WPr@  G?hA/.��X   WDTrA  G?nQz��;OX   PRPrB  G?XA/.��X   DTrC  G?b0�cV�X   ''rD  G?hA/.��X   PRP$rE  G?XA/.��X   JJSrF  G?XA/.��uhMjj  �rG  h h(h
c__builtin__
__main__
hNN}rH  NtrI  RrJ  �rK  RrL  (h�G?�[���\X   WRBrM  G?x��0�hMG?��a��X   INrN  G?��A)��X   NNrO  G?�z�ש{X   VBDrP  G?���|X   WPrQ  G?x��0�X   VBZrR  G?���|X   VBrS  G?x��0�X   TOrT  G?��A)��X   CCrU  G?���[��X   NNSrV  G?�`1�`X   VBNrW  G?x��0�X   CDrX  G?��A)��X   VBGrY  G?��A)��X   JJrZ  G?��A)��X   NNPr[  G?��A)��X   MDr\  G?x��0�X   POSr]  G?x��0�X   ``r^  G?x��0�uh�jL	  �r_  h h(h
c__builtin__
__main__
hNN}r`  Ntra  Rrb  �rc  Rrd  (X   JJre  G?�n2�e��X   NNrf  G?�t��y��X   RBSrg  G?�p"�E��X   NNPrh  G?�.\�X   NNSri  G?�h$�I��X   VBGrj  G?w@.�] �X   NNPSrk  G?� > | �X   ``rl  G?�p"�E��X   VBNrm  G?w@.�] �X   VBPrn  G?g@.�] �X   DTro  G?{ 6@l��X   JJSrp  G?� > | �X   VBDrq  G?s`&�M��X   RBrr  G?o > | �X   CDrs  G?�02`d��X   VBZrt  G?g@.�] �X   POSru  G?_ > | �X   JJRrv  G?s`&�M��h�G?o > | �X   INrw  G?o > | �X   WPrx  G?_ > | �X   VBry  G?_ > | �uX   INrz  j�  �r{  h h(h
c__builtin__
__main__
hNN}r|  Ntr}  Rr~  �r  Rr�  (X   NNPr�  G?�&L�2d�X   NNr�  G?�4hѣF�X   NNSr�  G?ͻv�۷oX   VBNr�  G?�(P�B�
X   INr�  G?�$H�"D�X   CDr�  G?�&L�2d�X   JJr�  G?ūV�Z�kX   WPr�  G?�0`��X   RBr�  G?� @�X   WRBr�  G?�0`��hMG?� @�X   VBGr�  G?�0`��X   DTr�  G?�0`��X   oovr�  G?� @�X   PRPr�  G?� @�X   VBPr�  G?�0`��X   VBr�  G?� @�X   VBZr�  G?� @�X   VBDr�  G?� @�uj�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   CCr�  G?�a�a�X   NNSr�  G?��0�1X   NNPr�  G?�UUUUUUX   NNPSr�  G?�a�a�X   NNr�  G?�I$�I$�X   JJr�  G?�a�a�h�G?�y�y�X   INr�  G?�y�y�X   WDTr�  G?�a�a�X   VBZr�  G?�a�a�X   POSr�  G?�a�a�X   VBDr�  G?�a�a�X   VBGr�  G?�a�a�uX   NNr�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   DTr�  G?�{�)���X   NNPr�  G?͞!��FX   VBr�  G?����^B�X   JJr�  G?�Pބ�@X   NNr�  G?��];<C�X   RBr�  G?��V��X   oovr�  G?�{�)���X   PRP$r�  G?p{�)���X   PRPr�  G?����'%�X   INr�  G?����}�X   NNSr�  G?����'%�X   TOr�  G?x�n��`RX   VBDr�  G?�{�)���X   VBNr�  G?p{�)���X   WRBr�  G?x�n��`RX   VBGr�  G?��n��`RX   VBZr�  G?��V��X   CDr�  G?��V��h�G?�Aj����X   JJRr�  G?p{�)���uj�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   NNPr�  G?�쎕3�X   NNr�  G?о�v�X   JJSr�  G?�H_
�;X   JJr�  G?���v�X   RBSr�  G?�쎕3�X   VBZr�  G?�쎕3�X   NNPSr�  G?�쎕3�X   ''r�  G?�쎕3�X   RBr�  G?�H_
�;X   NNSr�  G?�쎕3�X   CDr�  G?�H_
�;X   oovr�  G?�H_
�;X   VBGr�  G?�쎕3�X   DTr�  G?�H_
�;X   ``r�  G?�H_
�;uh�j1  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (NG?�+�+�X   VBNr�  G?�A�A�h�G?�A�A�X   INr�  G?�A�A�uj1  N�r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  NG?�      sNh%�r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   NNr�  G?׽����X   JJr�  G?�)�u�"�X   NNPr�  G?���9X   CDr�  G?�Ti*�GX   INr�  G?zJ�mQ��X   VBDr�  G?`���A	�X   RBSr�  G?s_{(!5�X   NNSr�  G?�����KX   JJSr�  G?�qxc��X   VBZr�  G?p���A	�X   JJRr�  G?q�;���X   NNPSr�  G?����A
X   ``r�  G?k�����X   VBNr�  G?`���A	�X   VBGr�  G?q�;���X   oovr�  G?`���A	�X   RBr�  G?`���A	�X   PRPr�  G?F#�wb@X   DTr�  G?P���A	�X   WDTr�  G?F#�wb@X   CCr�  G?P���A	�X   WPr�  G?F#�wb@uhMj'  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr   Rr  �r  Rr  (X   VBGr  G?��L�x��X   DTr  G?� ^)2�X   NNPr  G?ę�I�/X   NNr  G?�lߡ���X   VBr  G?���a{�X   PRPr	  G?���I�/X   JJr
  G?���a{�X   INr  G?���I�/X   NNSr  G?�lߡ���X   VBDr  G?��L�x��X   VBPr  G?��L�x��X   WPr  G?�lߡ���X   RBr  G?��L�x��X   CCr  G?���a{�X   PRP$r  G?��L�x��X   WRBr  G?��L�x��uj'  j  �r  h h(h
c__builtin__
__main__
hNN}r  Ntr  Rr  �r  Rr  (X   NNr  G?�q�q�X   DTr  G?�q�q�X   NNPr  G?�q�q�X   RPr  G?�UUUUUUX   ''r  G?�UUUUUUX   NNSr  G?�q�q�X   INr   G?�q�q�X   VBNr!  G?�q�q�X   ``r"  G?�UUUUUUX   TOr#  G?�q�q�uj  jX
  �r$  h h(h
c__builtin__
__main__
hNN}r%  Ntr&  Rr'  �r(  Rr)  (X   VBDr*  G?�ؼw\��h�G?��m�Kb�X   NNr+  G?����2A�X   INr,  G?��o�[�X   VBNr-  G?�a_;	lX   VBZr.  G?��*g��X   MDr/  G?�������X   NNSr0  G?�F�¿�|X   TOr1  G?�E�
�nX   VBPr2  G?�ؼw\��X   DTr3  G?�F�¿�|X   VBr4  G?�i:E�X   CCr5  G?�ؼw\��X   WRBr6  G?i �I��)X   JJr7  G?y �I��)X   RBr8  G?�ؼw\��X   oovr9  G?i �I��)X   WDTr:  G?�������X   VBGr;  G?i:E�hMG?� �I��)X   NNPr<  G?y �I��)X   RBSr=  G?i �I��)X   ``r>  G?i �I��)X   WPr?  G?i �I��)NG?y �I��)ujX
  j*  �r@  h h(h
c__builtin__
__main__
hNN}rA  NtrB  RrC  �rD  RrE  (X   VBNrF  G?�=�ҢX   WDTrG  G?�쎕3�X   RBrH  G?����n-^X   INrI  G?�Ң{#�X   NNPrJ  G?����n-^X   TOrK  G?�qj��&�X   DTrL  G?�* g�:TX   JJrM  G?�쎕3�X   oovrN  G?�qj��&�X   NNSrO  G?�qj��&�X   NNrP  G?�쎕3�h�G?�쎕3�uX   CDrQ  jX  �rR  h h(h
c__builtin__
__main__
hNN}rS  NtrT  RrU  �rV  RrW  (X   NNPrX  G?�uG�ƾX   POSrY  G?��uG�h�G?�Y9���}X   CDrZ  G?�!��>X   NNr[  G?�٤F��X   NNPSr\  G?�;��]�X   CCr]  G?�Y9���}X   VBDr^  G?�<�RF��X   JJr_  G?��uG�X   NNSr`  G?�洬U�~X   WDTra  G?j�/���X   TOrb  G?z�/���hMG?���E}X   INrc  G?�uG�ƾX   VBNrd  G?�U���X   ''re  G?a�uG�X   VBZrf  G?�U���X   RBrg  G?�U���X   VBrh  G?��r=��~X   VBPri  G?j�/���X   oovrj  G?q�uG�X   WPrk  G?v<�RF��X   MDrl  G?a�uG�ujd  h��rm  h h(h
c__builtin__
__main__
hNN}rn  Ntro  Rrp  �rq  Rrr  NG?�      shMj(  �rs  h h(h
c__builtin__
__main__
hNN}rt  Ntru  Rrv  �rw  Rrx  (X   NNPry  G?��؄u,�X   PRP$rz  G?�`���ϚX   NNr{  G?�ԲN��X   INr|  G?�K$�qZnX   WDTr}  G?��1��gX   TOr~  G?�1��g*X   DTr  G?��1��gX   CCr�  G?���@�X   WPr�  G?�`���ϚX   PRPr�  G?�ԲN��X   VBNr�  G?��1��ghMG?�ԲN��X   CDr�  G?��1��gX   NNSr�  G?��1��gh�G?�`���ϚX   JJr�  G?�x���C�X   MDr�  G?�`���ϚX   VBGr�  G?��1��gX   RPr�  G?�`���ϚX   JJSr�  G?�`���ϚX   oovr�  G?�`���ϚuX   VBNr�  h��r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (NG?��!k�X   NNr�  G?:�;��Dh�G?S�C��3X   ''r�  G?C�C��3X   ``r�  G?:�;��DX   NNPr�  G?:�;��DuX   NNPr�  h��r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   DTr�  G?���W���X   NNPr�  G?�`�vO��X   INr�  G?�9��q6X   RBr�  G?�zc���X   NNr�  G?�
2���X   TOr�  G?�`�vO��X   PRP$r�  G?�zc���X   VBNr�  G?���r;'�X   VBr�  G?����X   WRBr�  G?���𳁈X   NNSr�  G?�e���h�G?�zc���X   JJr�  G?���𳁈X   VBDr�  G?����X   WPr�  G?����X   VBZr�  G?pQ���4X   VBGr�  G?�e���X   oovr�  G?pQ���4X   JJSr�  G?pQ���4X   VBPr�  G?xzc���X   RPr�  G?xzc���X   PRPr�  G?����NG?pQ���4X   ''r�  G?pQ���4X   CDr�  G?xzc���uh�j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   NNr�  G?ނ�^���X   NNPr�  G?Ĺ��U	nX   JJr�  G?͞ݪ@fyX   JJSr�  G?�TSB X   VBNr�  G?y�'~|�X   VBGr�  G?v�xpo�X   CDr�  G?�1��u��X   VBZr�  G?qTSB X   NNSr�  G?���VvX   ``r�  G?qTSB X   oovr�  G?f�xpo�h�G?aTSB X   NNPSr�  G?���ba"VX   RBr�  G?f�xpo�X   INr�  G?s��ba"VX   JJRr�  G?qTSB X   DTr�  G?s��ba"VX   RBSr�  G?s��ba"VX   TOr�  G?V�xpo�X   VBDr�  G?V�xpo�X   CCr�  G?V�xpo�uX   INr�  j   �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   DTr�  G?�Jy��JX   JJr�  G?��cHzYX   PRPr�  G?��D}X   NNr�  G?��
���^X   RBr�  G?��A)��X   NNPr�  G?˘E';-�X   CDr�  G?�G%滂�X   VBPr�  G?uG%滂�X   NNSr�  G?���E';.X   INr�  G?�I��xZnX   oovr�  G?uG%滂�X   VBr�  G?���`jc�X   ''r�  G?uG%滂�X   PRP$r�  G?��D}X   VBGr�  G?uG%滂�X   JJSr�  G?uG%滂�X   NNPSr�  G?��D}X   JJRr�  G?�G%滂�X   VBNr�  G?uG%滂�X   TOr�  G?uG%滂�h�G?�A�A�uX   ''r�  j+  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (h�G?����u:X   INr�  G?ʸu9�7*X   NNr�  G?���HgoX   VBDr�  G?���Hgo1X   TOr�  G?���HgoX   ''r�  G?��֠R�[X   NNSr�  G?��+�#X   PRPr�  G?{�+�#X   VBZr�  G?��+�#X   VBr�  G?��+�#X   NNPr�  G?{�+�#X   VBNr�  G?�=2��vX   WRBr�  G?{�+�#X   DTr�  G?��+�#X   RBr�  G?��֠R�[X   WDTr�  G?{�+�#hMG?��֠R�[X   CCr   G?{�+�#X   VBGr  G?��+�#X   VBPr  G?��+�#X   MDr  G?{�+�#uX   VBDr  j�  �r  h h(h
c__builtin__
__main__
hNN}r  Ntr  Rr  �r	  Rr
  (X   VBNr  G?��7���h�G?����z�X   INr  G?ĺf�X[�X   JJr  G?����X   DTr  G?��ʾy
X   CCr  G?z���z�X   VBGr  G?���>�X   CDr  G?�5A����X   RBr  G?����E�X   NNPr  G?�Ɉ+�WX   VBr  G?����eX   TOr  G?���>�X   NNSr  G?����E�X   WPr  G?uɈ+�WhMG?x5A����X   oovr  G?c]�_�*�X   VBPr  G?c]�_�*�X   VBDr  G?m��n�tX   JJRr  G?s]�_�*�X   NNr  G?�W& �LAX   WRBr  G?m��n�tX   VBZr  G?h5A����X   ``r  G?]��n�tX   PRPr   G?S]�_�*�X   NNPSr!  G?]��n�tX   WDTr"  G?S]�_�*�uj�  j  �r#  h h(h
c__builtin__
__main__
hNN}r$  Ntr%  Rr&  �r'  Rr(  (h�G?�=H'�c�X   INr)  G?޻��1�X   TOr*  G?�K�D�kX   JJSr+  G?G �GA�X   NNr,  G?����{�X   WRBr-  G?|���X   JJr.  G?�ı�A<KX   NNSr/  G?����*${X   RPr0  G?{P�ؤ��X   VBNr1  G?�4�ڵ�cX   ''r2  G?i���0)�X   DTr3  G?�,��X   VBDr4  G?Q@�Euq!X   WPr5  G?�p�����X   VBGr6  G?w �GA�X   CCr7  G?����;7X   JJRr8  G?Q@�Euq!X   PRP$r9  G?a@�Euq!X   RBr:  G?�P�ؤ��X   PRPr;  G?a@�Euq!X   NNPr<  G?�y	ASK�hMG?t �&^YQX   oovr=  G?g �GA�X   ``r>  G?a@�Euq!X   WDTr?  G?Q@�Euq!X   MDr@  G?G �GA�NG?W �GA�X   CDrA  G?G �GA�X   VBZrB  G?G �GA�ujg  h��rC  h h(h
c__builtin__
__main__
hNN}rD  NtrE  RrF  �rG  RrH  NG?�      sX   JJrI  jx  �rJ  h h(h
c__builtin__
__main__
hNN}rK  NtrL  RrM  �rN  RrO  (X   NNrP  G?�s#:�X   VBNrQ  G?�.��A��X   INrR  G?�#:�1R4X   JJrS  G?�|z �w�X   NNPSrT  G?���M�,�h�G?���M�,�X   VBGrU  G?���M�,�X   VBrV  G?���M�,�X   NNSrW  G?���M�,�X   NNPrX  G?���M�,�X   RBrY  G?���M�,�ujx  jP  �rZ  h h(h
c__builtin__
__main__
hNN}r[  Ntr\  Rr]  �r^  Rr_  (X   VBDr`  G?����.�X   POSra  G?at]E�tX   NNrb  G?�E�t]X   CDrc  G?gE�t]FX   PRPrd  G?mE�t]X   INre  G?�.���/X   JJrf  G?z.���/X   VBNrg  G?�.���/h�G?���.��X   NNSrh  G?��.���hMG?��.���X   VBGri  G?}E�t]X   TOrj  G?�E�t]X   NNPrk  G?�t]E�tX   RBrl  G?��.���X   VBZrm  G?}E�t]X   WDTrn  G?z.���/X   DTro  G?��t]E�X   ''rp  G?qt]E�tX   CCrq  G?qt]E�tX   VBPrr  G?WE�t]FX   VBrs  G?gE�t]FX   WRBrt  G?at]E�tNG?WE�t]FX   oovru  G?at]E�tX   ``rv  G?WE�t]FuNh&�rw  h h(h
c__builtin__
__main__
hNN}rx  Ntry  Rrz  �r{  Rr|  (X   NNPr}  G?��o��o�X   DTr~  G?��o��o�X   NNr  G?͉؝�؞X   PRPr�  G?�A�A�X   INr�  G?��;�;X   VBr�  G?�A�A�X   NNSr�  G?��;�;X   JJr�  G?�A�A�X   WRBr�  G?�A�A�X   oovr�  G?�A�A�uh&j}  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   POSr�  G?���F~%X   ''r�  G?���J3�X   NNPSr�  G?}�`v���X   INr�  G?���J3�X   NNPr�  G?��k��X   VBZr�  G?�g�Q��FX   NNr�  G?��`v���X   DTr�  G?}�`v���h�G?�B�Y!dX   CCr�  G?���g�Q�X   TOr�  G?��`v���X   PRPr�  G?���J3�)X   CDr�  G?m�`v���X   NNSr�  G?��`v���X   JJr�  G?}�`v���X   oovr�  G?�B�Y!dX   VBDr�  G?vB�Y!dhMG?���J3�)X   ``r�  G?���J3�)X   RBr�  G?vB�Y!dX   VBr�  G?vB�Y!duj�  jP  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   ''r�  G?�UUUUUUX   VBNr�  G?�UUUUUUX   NNr�  G?�UUUUUUujP  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   VBDr�  G?�򆼡�(h�G?�C^Pה6X   NNr�  G?�5�yC^X   VBPr�  G?�򆼡�(X   TOr�  G?�򆼡�(NG?�5�yC^X   INr�  G?�5�yC^X   VBNr�  G?�򆼡�(uj�  jG  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   JJr�  G?�      X   NNr�  G?�      X   CDr�  G?�X   INr�  G?�X   MDr�  G?�������X   VBDr�  G?�UUUUUUX   JJSr�  G?�X   VBZr�  G?�������X   VBPr�  G?�X   NNSr�  G?�UUUUUUX   RBr�  G?�X   VBGr�  G?�X   NNPr�  G?�uj�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   DTr�  G?���n/N�X   PRP$r�  G?�����J�X   INr�  G?��x�]�X   NNPr�  G?�G�k}tyX   NNr�  G?�vDݑ7X   CCr�  G?L�m���h�G?����i�X   WPr�  G?�)�d2�X   JJRr�  G?jY9Ɂ��X   JJr�  G?�tŝ1gLX   VBGr�  G?�]����X   NNSr�  G?���i���X   PRPr�  G?��l�lX   CDr�  G?��б@�X   JJSr�  G?q�}�pX   WDTr�  G?t\8JAE�X   oovr�  G?e��0�X�X   VBNr�  G?e��0�X�X   WRBr�  G?e��0�X�X   RBr�  G?s)�d2�X   ``r�  G?jY9Ɂ��hMG?S)�d2�X   NNPSr�  G?C)�d2�NG?S)�d2�X   TOr�  G?L�m���X   VBDr�  G?S)�d2�X   POSr�  G?C)�d2�X   VBZr�  G?C)�d2�uX   NNr�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (h�G?��i�!�X   INr�  G?ƹ��n,TX   NNr�  G?��(x�ܫX   VBNr�  G?�<b�Up�X   NNPr�  G?��y qX   VBZr�  G?�E�����X   TOr�  G?�����1X   RBr�  G?� qa�lX   PRPr�  G?cE�����hMG?�`
GN��X   VBDr�  G?���6H�X   VBPr�  G?�Ӭ|��.X   WDTr�  G?�3O,�X   DTr�  G?�<b�Up�X   ''r�  G?g qa�lX   VBGr�  G?�E�����X   JJr�  G?����t��X   MDr�  G?� qa�lX   oovr�  G?lDiZ�X   RPr�  G?W qa�lX   CCr   G?����t��X   NNSr  G?t��c��X   VBr  G?��6��XX   CDr  G?T��c��X   WPr  G?n��ׇ:X   WRBr  G?q�ɷhd7X   RBSr  G?I�D��FX   POSr  G?d��c��X   JJRr  G?I�D��FNG?g qa�lX   ``r	  G?I�D��FX   PRP$r
  G?I�D��FX   NNPSr  G?4��c��uj5  j�  �r  h h(h
c__builtin__
__main__
hNN}r  Ntr  Rr  �r  Rr  (X   JJr  G?��=���X   NNPr  G?�{���aX   DTr  G?���a|X   NNSr  G?��i�XGX   PRPr  G?���a|X   VBNr  G?���a{�X   NNr  G?Ѝ=���X   VBr  G?���a{�X   CDr  G?���a|X   oovr  G?�{���aX   NNPSr  G?���a{�h�G?�{���aX   INr  G?���a|X   VBZr  G?���a{�X   TOr  G?�{���aX   VBGr   G?���a{�X   RBr!  G?���a{�uj�  j  �r"  h h(h
c__builtin__
__main__
hNN}r#  Ntr$  Rr%  �r&  Rr'  (X   NNPr(  G?�
b�H-�X   ''r)  G?��� 1�X   CDr*  G?� ���5|X   NNr+  G?��I�~��X   INr,  G?x��zEX   JJr-  G?���zEX   NNSr.  G?�,�>O��X   VBGr/  G?x��zEhMG?����s�X   TOr0  G?p�ۦ��`h�G?��ۦ��`X   NNPSr1  G?� ���5|X   CCr2  G?��R�[d8X   ``r3  G?���zEX   VBZr4  G?p�ۦ��`X   MDr5  G?p�ۦ��`uX   NNPr6  j	  �r7  h h(h
c__builtin__
__main__
hNN}r8  Ntr9  Rr:  �r;  Rr<  (X   ''r=  G?���X   VBDr>  G?�SgSgX   VBPr?  G?ǿ!��!�h�G?Ё�Ё��X   VBZr@  G?�����X   INrA  G?�*�*�hMG?�����X   WRBrB  G?�����X   NNSrC  G?���X   NNPSrD  G?�����X   DTrE  G?�*�*�X   POSrF  G?���X   NNPrG  G?�����X   CCrH  G?�*�*�X   NNrI  G?�7�7�X   RBrJ  G?���X   VBrK  G?�7�7�X   JJrL  G?�����X   MDrM  G?���X   TOrN  G?���uj	  j=  �rO  h h(h
c__builtin__
__main__
hNN}rP  NtrQ  RrR  �rS  RrT  (X   NNrU  G?�      X   VBDrV  G?�UUUUUUh�G?ڪ�����X   NNSrW  G?�UUUUUUuNh'�rX  h h(h
c__builtin__
__main__
hNN}rY  NtrZ  Rr[  �r\  Rr]  (X   JJr^  G?�UUUUUUX   NNr_  G?��8�9X   NNSr`  G?�UUUUUUX   JJSra  G?�q�q�uhMj)  �rb  h h(h
c__builtin__
__main__
hNN}rc  Ntrd  Rre  �rf  Rrg  (hMG?�nF�nF�h�G?�V�jV�jX   INrh  G?���؝��X   NNPri  G?��nF�nGX   VBDrj  G?�jV�jV�X   RBrk  G?��;�;X   POSrl  G?��;�;X   oovrm  G?w�z�zX   CCrn  G?�ннX   CDro  G?��؝�؞X   VBNrp  G?s�;�;X   VBPrq  G?�����X   VBZrr  G?��z�zX   NNrs  G?��؝�؞X   NNSrt  G?{����X   VBru  G?g�z�zX   MDrv  G?g�z�zX   DTrw  G?_���� X   NNPSrx  G?���� X   PRPry  G?_���� X   WPrz  G?_���� X   JJr{  G?g�z�zX   TOr|  G?o���� X   ``r}  G?o���� uX   VBDr~  j�	  �r  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   JJr�  G?�r��8h�G?���G��X   PRPr�  G?�[�
��X   NNPr�  G?���w��X   DTr�  G?���G��X   NNSr�  G?�M"���X   CDr�  G?��f�ߔ�X   NNr�  G?�M"����X   RBr�  G?��f�ߔ�X   JJRr�  G?���;?�tX   VBZr�  G?���;?�tX   VBNr�  G?���;?�tX   VBGr�  G?��f�ߔ�X   NNPSr�  G?���;?�tX   TOr�  G?���;?�tX   WRBr�  G?���;?�tX   WPr�  G?���;?�tX   PRP$r�  G?���;?�tX   MDr�  G?���;?�tX   oovr�  G?���;?�tuj�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   INr�  G?�T�ۖ�h�G?��ۖ��X   JJr�  G?���<�LX   NNr�  G?�탤!�JX   VBDr�  G?�?�&�X   VBNr�  G?�Ibת�X   VBZr�  G?����/�iX   TOr�  G?z�nZ��rX   CCr�  G?��$����X   RBr�  G?�*���VX   WDTr�  G?z�nZ��rX   VBr�  G?��nZ��rX   NNPSr�  G?q��<�LX   DTr�  G?q��<�LX   NNSr�  G?���<�LX   ``r�  G?z�nZ��rX   VBPr�  G?z�nZ��rNG?�h1K��_X   VBGr�  G?�h1K��_hMG?�h1K��_X   MDr�  G?���<�LX   oovr�  G?���<�LX   NNPr�  G?���<�LX   ''r�  G?q��<�Luj�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   DTr�  G?�,��,X   WDTr�  G?��!B�X   CDr�  G?��9�s��h�G?�D�4MEX   NNPr�  G?���?O��X   JJr�  G?��`XX   NNr�  G?��yG��X   NNSr�  G?��`XX   VBGr�  G?��`XX   WPr�  G?��!B�X   POSr�  G?��`XX   PRP$r�  G?��1�c�X   INr�  G?�D�4MEX   PRPr�  G?�D�4MEX   ``r�  G?��`XuX   VBr�  j  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   INr�  G?۔�Y��h�G?�k�r.��X   NNPr�  G?�G}�)"X   VBNr�  G?�"}�Q��X   TOr�  G?��mx.FX   VBGr�  G?����lX   DTr�  G?�Ǩ��dX   PRP$r�  G?d����X   NNSr�  G?��cf�=�X   JJr�  G?��<2���X   RPr�  G?�#X�]03X   NNr�  G?������X   RBr�  G?��۔�ZX   WPr�  G?}"}�Q��X   WRBr�  G?��s
�hMG?t����X   oovr�  G?d����X   VBr�  G?[k�r.��X   ``r�  G?[k�r.��X   CCr�  G?}"}�Q��X   VBPr�  G?T����X   WDTr�  G?Kk�r.��X   JJRr�  G?kk�r.��X   PRPr�  G?Kk�r.��X   CDr�  G?a#X�]03NG?Kk�r.��X   NNPSr�  G?Kk�r.��X   ''r�  G?Kk�r.��X   VBZr�  G?T����X   VBDr�  G?Kk�r.��uj�  j-  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   NNr�  G?���'12�X   NNSr�  G?�qh<
h�G?�U���X   VBDr�  G?�Y9���}X   NNPr�  G?�Xd�r>X   JJr�  G?�� �k��X   INr�  G?�Y9���}X   VBZr�  G?��r=��~X   VBGr�  G?z�/���X   NNPSr�  G?z�/���X   RBr�  G?z�/���X   ``r�  G?z�/���uj  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   INr   G?����+c�X   ''r  G?���+c��X   NNr  G?�<��N	h�G?���/��X   CCr  G?�I�A��X   NNPr  G?�����8hX   TOr  G?���+c��X   MDr  G?��I�A�hMG?��Ely}�X   VBZr  G?����8h#X   VBNr  G?�p�Ely~X   POSr	  G?�4[_uX   RBr
  G?�[_u'X   VBDr  G?�A���RX   VBPr  G?��A���X   CDr  G?a[_u'X   VBr  G?���+c��X   VBGr  G?�[_u'NG?j��/��X   JJr  G?���+c��X   NNSr  G?�p�Ely~X   NNPSr  G?u���Rp�X   WPr  G?~_u'WX   DTr  G?j��/��X   WDTr  G?j��/��X   WRBr  G?a[_u'uj�  j   �r  h h(h
c__builtin__
__main__
hNN}r  Ntr  Rr  �r  Rr  (X   NNPr  G?��~��X   WPr  G?�n5ͪ�X   CDr  G?��~��X   DTr   G?���;�xX   NNr!  G?���e�>{X   WDTr"  G?�[_u'X   INr#  G?�=�9FKX   NNPSr$  G?�Ӿ&.�X   RBr%  G?{��e�>{X   PRP$r&  G?���~��h�G?���e�>{X   ``r'  G?�Ӿ&.�X   VBGr(  G?���e�>{X   NNSr)  G?���e�>{X   VBZr*  G?{��e�>{X   JJr+  G?�[_u'X   TOr,  G?�Ӿ&.�X   WRBr-  G?{��e�>{X   PRPr.  G?{��e�>{uj�  j�  �r/  h h(h
c__builtin__
__main__
hNN}r0  Ntr1  Rr2  �r3  Rr4  (X   PRPr5  G?�.��A��X   ''r6  G?�|z �w�X   INr7  G?�p���X   DTr8  G?��8]��X   RBr9  G?�.��A��X   VBNr:  G?�.��A��hMG?���M�,�X   NNPr;  G?�.��A��X   NNr<  G?�|z �w�X   JJr=  G?�|z �w�h�G?�|z �w�X   TOr>  G?�.��A��X   CDr?  G?���M�,�X   POSr@  G?���M�,�X   ``rA  G?�չ���\X   RPrB  G?���M�,�X   PRP$rC  G?���M�,�uj5  j  �rD  h h(h
c__builtin__
__main__
hNN}rE  NtrF  RrG  �rH  RrI  (X   ''rJ  G?�q�q�h�G?�UUUUUUX   INrK  G?�q�q�X   NNSrL  G?�q�q�X   TOrM  G?�q�q�X   DTrN  G?�q�q�uj  jJ  �rO  h h(h
c__builtin__
__main__
hNN}rP  NtrQ  RrR  �rS  RrT  (X   RBrU  G?�      X   NNrV  G?�      X   NNSrW  G?�      ujJ  jU  �rX  h h(h
c__builtin__
__main__
hNN}rY  NtrZ  Rr[  �r\  Rr]  (X   JJr^  G?�������X   VBNr_  G?�\(��X   INr`  G?�(�\)X   VBZra  G?��Q��X   VBPrb  G?�z�G�{X   VBDrc  G?�z�G�{X   VBrd  G?�z�G�{X   RBre  G?�z�G�{ujU  j^  �rf  h h(h
c__builtin__
__main__
hNN}rg  Ntrh  Rri  �rj  Rrk  (X   NNrl  G?��ǧ�:X   INrm  G?�s#��h�G?��SJ��hX   CCrn  G?��~�+GtX   NNSro  G?�Ò��_"X   RBrp  G?�c7�<X   TOrq  G?��0-��X   JJrr  G?�;3�o�VhMG?�%���owX   NNPrs  G?��~�+GtX   PRPrt  G?j!z�u�/X   MDru  G?c�,cX   WPrv  G?pT��i�}X   ''rw  G?v�K��?IX   VBNrx  G?s�,cX   JJRry  G?Z!z�u�/X   WRBrz  G?z!z�u�/X   VBGr{  G?}e�B$�X   WDTr|  G?c�,cX   VBPr}  G?c�,cX   PRP$r~  G?Z!z�u�/X   oovr  G?c�,cX   CDr�  G?c�,cNG?j!z�u�/X   DTr�  G?c�,cX   VBZr�  G?c�,cX   NNPSr�  G?Z!z�u�/X   VBDr�  G?Z!z�u�/X   ``r�  G?c�,cuX   INr�  jL  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   NNr�  G?ب�����X   NNSr�  G?�<�<�h�G?��@�@X   CDr�  G?s�8�8X   CCr�  G?�X   VBGr�  G?}A�A�X   TOr�  G?r[�[�X   JJr�  G?�G"�G"�X   NNPr�  G?�����X   INr�  G?�Y~Y~X   VBDr�  G?n�h�hX   NNPSr�  G?�D�D hMG?w�<�<X   VBNr�  G?n�h�hX   WPr�  G?T����X   WDTr�  G?2[�[�X   MDr�  G?B[�[�X   VBPr�  G?l����X   VBZr�  G?d����X   ``r�  G?B[�[�X   DTr�  G?F�`�`X   VBr�  G?T����X   WRBr�  G?V�`�`X   JJRr�  G?;�@�@X   RBr�  G?Y=�=�X   oovr�  G?PNG?F�`�`X   RBSr�  G?2[�[�X   PRPr�  G?2[�[�X   JJSr�  G?2[�[�X   RPr�  G?2[�[�X   POSr�  G?;�@�@uj�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   INr�  G?�З�%�	X   JJr�  G?�q�q�X   ``r�  G?���%�	{X   DTr�  G?͡/hK�X   NNr�  G?�З�%�	X   RBr�  G?�UUUUUUX   VBNr�  G?�����/hX   VBDr�  G?�q�q�X   NNPr�  G?���%�	{X   CDr�  G?�З�%�	X   VBZr�  G?�q�q�X   NNSr�  G?�����/hX   CCr�  G?�����/hh�G?�����/hX   PRPr�  G?�����/hX   VBGr�  G?�����/huj�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   DTr�  G?��vr�X   WPr�  G?���@�X   RBr�  G?���@�X   NNSr�  G?�1��g*X   JJr�  G?��vr�zh�G?��1��gX   NNr�  G?��1��gX   NNPr�  G?��1��gX   INr�  G?��1��gX   PRPr�  G?��vr�X   PRP$r�  G?���@�X   JJRr�  G?��1��gX   JJSr�  G?��1��gX   CDr�  G?���@�X   VBr�  G?��1��gX   VBNr�  G?��1��guX   ''r�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (h�G?�I$�I$�X   NNr�  G?ݶ�m��nX   INr�  G?�m��m��X   NNSr�  G?�m��m��X   VBDr�  G?�I$�I$�X   CDr�  G?�m��m��uj�  j  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   DTr�  G?��L�oj�X   INr�  G?�Rńu�aX   NNPr�  G?�Ĝ��ͨX   PRPr�  G?���:f�X   VBNr�  G?���h��h�G?�
�[\nX   VBDr�  G?o�6�	
�X   JJr�  G?�P�B��X   WPr�  G?��/���PX   JJRr�  G?{�/���PX   RBr�  G?�{�,��X   NNSr�  G?�Fq/#��X   TOr�  G?�����zdX   JJSr�  G?biu+���X   WRBr�  G?x����}�X   NNr�  G?��)�RqYX   PRP$r�  G?�?_��:'X   VBGr�  G?�?_��:'X   CDr�  G?riu+���X   RPr�  G?�Ĝ��ͨX   NNPSr�  G?W�(���X   VBr�  G?o�6�	
�X   CCr�  G?jM�в3�X   oovr�  G?sˤ��X   VBZr�  G?n?��3T�hMG?a�:�;X   WDTr�  G?ZM�в3�X   VBPr�  G?_�6�	
�X   ``r   G?W�(���X   RBSr  G?g�(���X   MDr  G?\�ܲ]�NG?_�6�	
�X   POSr  G?5
�[\nuX   DTr  j�  �r  h h(h
c__builtin__
__main__
hNN}r  Ntr  Rr  �r	  Rr
  (X   NNr  G?�x,!��PX   JJr  G?����6X   NNSr  G?�Ĩ�1�>X   VBGr  G?����6X   RBr  G?!� ��X   INr  G?����6X   NNPr  G?���5 �hMG?g���6X   PRPr  G?S�}�6�X   VBNr  G?���5 �h�G?�K���AtX   VBDr  G?\�m�OQ�X   CCr  G?��D���)X   WPr  G?p�����X   TOr  G?g���6X   DTr  G?s�}�6�X   CDr  G?l�m�OQ�X   NNPSr  G?S�}�6�X   ``r  G?c�}�6�X   VBZr  G?S�}�6�X   JJSr  G?S�}�6�uj  j�	  �r  h h(h
c__builtin__
__main__
hNN}r  Ntr   Rr!  �r"  Rr#  (X   INr$  G?ބr��GX   TOr%  G?��ô�[�h�G?�.t���X   JJr&  G?����X   NNPr'  G?������X   RPr(  G?�ı�A<KX   RBr)  G?�ʠ��X   NNSr*  G?��ô�[�X   VBZr+  G?o���X   JJRr,  G?o���X   DTr-  G?��ô�[�X   CCr.  G?�ı�A<KX   VBGr/  G?w���{�X   NNr0  G?������X   VBNr1  G?��ô�[�hMG?����X   WPr2  G?w���{�X   VBr3  G?o���X   oovr4  G?���X   WRBr5  G?w���{�X   ``r6  G?o���NG?o���X   WDTr7  G?o���X   JJSr8  G?w���{�uX   VBNr9  j�  �r:  h h(h
c__builtin__
__main__
hNN}r;  Ntr<  Rr=  �r>  Rr?  (h�G?�v�Wj%wX   INr@  G?������X   VBPrA  G?������X   NNrB  G?�81�8X   WRBrC  G?��Q+��X   JJrD  G?�ډ]���X   VBZrE  G?������X   VBDrF  G?������X   RBrG  G?x�����X   TOrH  G?��Q+��X   PRPrI  G?x�����X   MDrJ  G?x�����X   oovrK  G?x�����X   CCrL  G?x�����uj�  h��rM  h h(h
c__builtin__
__main__
hNN}rN  NtrO  RrP  �rQ  RrR  NG?�      sX   JJrS  jR  �rT  h h(h
c__builtin__
__main__
hNN}rU  NtrV  RrW  �rX  RrY  (X   ``rZ  G?|����MX   NNPr[  G?èn̟�X   PRPr\  G?���'�X   VBDr]  G?��n̟�X   NNr^  G?���'�X   DTr_  G?ڱФip$X   VBGr`  G?|����MX   JJra  G?�q�<PkX   VBZrb  G?��n̟�X   RBrc  G?��1%��X   NNSrd  G?�q�<Pk:X   INre  G?�;k��~X   VBNrf  G?��'�=5*X   oovrg  G?l����MX   WRBrh  G?uq�<Pk:X   VBPri  G?|����MX   JJSrj  G?|����MX   CDrk  G?���'�X   MDrl  G?l����MX   VBrm  G?���\�X   JJRrn  G?l����MX   WPro  G?���\�X   TOrp  G?uq�<Pk:X   RPrq  G?l����MX   RBSrr  G?l����MX   PRP$rs  G?|����MujR  jZ  �rt  h h(h
c__builtin__
__main__
hNN}ru  Ntrv  Rrw  �rx  Rry  (X   NNPrz  G?��~��~�X   DTr{  G?�-�-�X   JJr|  G?��~��~�X   CDr}  G?��h�hX   NNr~  G?��h�hX   VBr  G?���X   NNSr�  G?�!�!�X   VBGr�  G?��h�hX   INr�  G?��h�hX   RBr�  G?���X   PRP$r�  G?��h�hX   VBNr�  G?��h�hX   TOr�  G?��h�hh�G?��h�hX   CCr�  G?��h�hX   PRPr�  G?���ujS  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   NNSr�  G?Ӣ�-�f�X   CCr�  G?��5�x��X   JJr�  G?�ڷ��CX   NNPr�  G?�gd�oX   INr�  G?���W��X   NNr�  G?�!�L�h�G?�e�%H�hMG?��G��jX   TOr�  G?��5�x��X   VBZr�  G?�G��jX   ''r�  G?��>��X   VBDr�  G?��5�x��X   POSr�  G?��,��X   WPr�  G?o�G��jX   VBGr�  G?�G��jX   JJSr�  G?��(C��X   VBNr�  G?��(C��X   RBr�  G?w�5�x��X   CDr�  G?w�5�x��NG?w�5�x��X   ``r�  G?o�G��jujs  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   NNr�  G?�t�y��GX   INr�  G?�Tp�}X   NNSr�  G?� *��x�h�G?�Ͽ�8KX   VBDr�  G?� *��x�X   JJr�  G?�o>���,X   TOr�  G?� *��x�X   VBZr�  G?�|�2�oX   NNPr�  G?��h�d�X   CDr�  G?�ï��]�X   DTr�  G?uq�<Pk:X   VBGr�  G?��h�d�NG?uq�<Pk:X   RBr�  G?�ï��]�X   MDr�  G?�q�<PkX   VBr�  G?�q�<PkX   VBNr�  G?uq�<Pk:uj�  j?  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   TOr�  G?���6��X   oovr�  G?�i���HX   INr�  G?�Lo��X   JJSr�  G?}T��
�X   VBNr�  G?��A�?X   RBr�  G?��c|��X   JJr�  G?��A�?X   NNPr�  G?�i���HX   PRPr�  G?����H��X   DTr�  G?��#/QJh�G?���]k�&hMG?si���HX   WPr�  G?�T��
�X   VBGr�  G?�2��&�X   NNSr�  G?��#/QJX   PRP$r�  G?�i���HX   ''r�  G?�T��
�X   VBDr�  G?�C�pՉX   JJRr�  G?�T��
�X   NNr�  G?�X����X   VBr�  G?�i���HX   VBZr�  G?}T��
�X   WRBr�  G?si���HX   RBSr�  G?si���HX   RPr�  G?�C�pՉX   CDr�  G?�C�pՉX   VBPr�  G?si���HX   ``r�  G?�C�pՉuj?  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   PRPr�  G?p�Dc��X   DTr�  G?�'��Z�X   NNPr�  G?�K3����h�G?�'��Z�X   VBr�  G?�R��t�X   INr�  G?���¯�X   NNSr�  G?�@2O!�+X   WRBr�  G?i'��Z�X   NNr�  G?��N|vpX   PRP$r�  G?�ݬ��1X   JJr�  G?�@2O!�+X   RBr�  G?p�Dc��X   RBSr�  G?i'��Z�X   WPr�  G?�ݬ��1X   NNPSr�  G?`�Dc��X   WDTr�  G?`�Dc��X   VBGr�  G?}Xӷ�?iX   TOr�  G?`�Dc��X   JJRr�  G?`�Dc��X   CDr�  G?`�Dc��uj�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   ''r�  G?���k�h�G?�!�~u4oX   INr�  G?�M�P1YhMG?���ː��X   VBr�  G?���ː��X   VBZr�  G?���k�X   CCr�  G?���ː��X   VBGr�  G?���k�X   DTr�  G?���k�X   RBr�  G?���k�X   JJSr�  G?���k�X   TOr�  G?���k�X   WPr�  G?���k�uX   CDr   jY  �r  h h(h
c__builtin__
__main__
hNN}r  Ntr  Rr  �r  Rr  (X   NNPr  G?�X��Ƈ�X   NNSr  G?��_�_X   NNr	  G?�2�	G�X   CDr
  G?p���%��X   JJr  G?��1Ί��h�G?����%��X   TOr  G?����%��X   VBNr  G?p���%��X   INr  G?��+���X   CCr  G?vJ�:��_X   NNPSr  G?p���%��X   VBGr  G?��+���X   VBZr  G?fJ�:��_X   RBr  G?p���%��ujY  jQ  �r  h h(h
c__builtin__
__main__
hNN}r  Ntr  Rr  �r  Rr  (h�G?�*ً�V�X   VBPr  G?ų���X   VBDr  G?�0W塂�X   VBNr  G?���=�X   MDr  G?�+���_�X   TOr  G?�+���_�X   INr  G?� ���X   RBr   G?�Ò ��X   CCr!  G?�w�x۾X   WDTr"  G?q�S����X   VBZr#  G?�^}@���X   RBSr$  G?j^}@���X   POSr%  G?�Ò ��X   NNr&  G?�����l�hMG?����6�X   VBr'  G?�{H��rX   VBGr(  G?����6�X   oovr)  G?j^}@���X   PRPr*  G?q�S����X   NNSr+  G?u�h`��CX   CDr,  G?a�S����X   DTr-  G?j^}@���NG?j^}@���X   ''r.  G?a�S����X   WRBr/  G?q�S����X   JJr0  G?u�h`��CX   WPr1  G?a�S����uX   PRP$r2  j�  �r3  h h(h
c__builtin__
__main__
hNN}r4  Ntr5  Rr6  �r7  Rr8  (X   INr9  G?��vr�X   NNr:  G?�~��@�X   NNPr;  G?зg*�LX   JJSr<  G?��1��gX   CCr=  G?���@�h�G?���1��X   VBr>  G?��1��gX   POSr?  G?���@�X   NNSr@  G?��1��gX   TOrA  G?���@�X   VBNrB  G?��1��gX   VBZrC  G?���@�hMG?��1��gX   VBDrD  G?��1��gX   ``rE  G?���@�uX   NNPrF  js  �rG  h h(h
c__builtin__
__main__
hNN}rH  NtrI  RrJ  �rK  RrL  (X   VBrM  G?吲B�YX   NNSrN  G?yp���rX   RBrO  G?��֨��X   NNrP  G?��6�X   PRPrQ  G?���O�X   ``rR  G?yp���rX   CDrS  G?�p���rX   NNPrT  G?���	�Vh�G?�p���rX   TOrU  G?yp���rX   VBNrV  G?yp���rX   VBDrW  G?���	�VX   DTrX  G?�B�Y!dujs  jM  �rY  h h(h
c__builtin__
__main__
hNN}rZ  Ntr[  Rr\  �r]  Rr^  (X   INr_  G?��b/�X   VBDr`  G?xc��i��X   DTra  G?�b/�s9X   PRPrb  G?�<�]�ߊX   NNrc  G?���|wX   VBNrd  G?��@��X   NNPre  G?���ph�G?�ہc̵�X   NNSrf  G?�p,y��X   JJrg  G?��sf�-X   VBrh  G?�����X   POSri  G?d���5CX   VBGrj  G?����0�`X   RBrk  G?��W?	<X   JJRrl  G?~ �vsO�X   TOrm  G?��'���X   CDrn  G?v�n�'MX   WRBro  G?�<�]�ߊX   VBZrp  G?F�n�'MX   PRP$rq  G?������VX   WPrr  G?�#��+}X   CCrs  G?|���0�`X   RPrt  G?v�n�'MX   MDru  G?Q7SR:X   oovrv  G?d���5CX   VBPrw  G?F�n�'MX   WDTrx  G?d���5ChMG?\���0�`X   ``ry  G?a7SR:X   ''rz  G?Q7SR:X   RBSr{  G?f�n�'MX   JJSr|  G?Q7SR:uX   NNr}  j  �r~  h h(h
c__builtin__
__main__
hNN}r  Ntr�  Rr�  �r�  Rr�  (X   VBDr�  G?�����X   NNPr�  G?�r��pM�X   VBZr�  G?�.G�)��X   VBPr�  G?�/�A��4X   MDr�  G?�	b���PX   NNSr�  G?���/@g�X   NNr�  G?���ajzVX   RBr�  G?���,��~X   DTr�  G?r��!�xX   JJr�  G?�MY��X   CDr�  G?o��^өX   INr�  G?o��^өX   NNPSr�  G?T�����uj  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   INr�  G?�J��nX   NNr�  G?������X   PRPr�  G?�5�U� �X   VBNr�  G?��u �%X   NNPr�  G?���l��X   RBr�  G?���oU|X   JJr�  G?��PD�X   NNSr�  G?����|�X   TOr�  G?�M�[�R�X   DTr�  G?����0�X   VBGr�  G?�e[aF��X   JJRr�  G?�Sq��y�X   RPr�  G?�ėw�MRX   CDr�  G?}J��nX   PRP$r�  G?���l��h�G?eėw�MRX   WPr�  G?uėw�MRX   CCr�  G?uėw�MRhMG?]J��nX   RBSr�  G?eėw�MRX   oovr�  G?r#ӎ��X   VBr�  G?eėw�MRX   VBDr�  G?]J��nX   JJSr�  G?]J��nX   ``r�  G?eėw�MRX   WRBr�  G?eėw�MRuX   NNr�  j  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   PRPr�  G?���[��X   JJr�  G?�b@h�<�h�G?�b@h�<�X   INr�  G?��l�b�%X   NNPr�  G?�3O%���X   DTr�  G?Ǿ�!לX   VBDr�  G?�]�F�X   NNr�  G?�Fi�8X   RBr�  G?�3O%���X   VBNr�  G?�b@h�<�X   TOr�  G?�w�քX   NNSr�  G?��l�b�%X   MDr�  G?�3O%���X   WPr�  G?�w�քX   VBGr�  G?������X   CDr�  G?�3O%���X   VBZr�  G?�w�քX   NNPSr�  G?z3O%���X   ``r�  G?qw�քhMG?qw�քX   VBPr�  G?z3O%���X   PRP$r�  G?z3O%���X   JJSr�  G?z3O%���X   oovr�  G?�w�քX   WDTr�  G?qw�քuj@  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   ``r�  G?�X   JJr�  G?�X   INr�  G?ϟ�����X   TOr�  G?�X   DTr�  G?�X   ''r�  G?�h�G?ə�����X   VBDr�  G?�X   MDr�  G?�hMG?�X   NNr�  G?�X   NNSr�  G?�X   RBr�  G?�X   NNPr�  G?�X   CCr�  G?�X   VBr�  G?�X   JJRr�  G?�uj�  j)  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   VBr�  G?�����X   INr�  G?�F�F�h�G?�7�7�X   VBZr�  G?���X   VBNr�  G?�7�7�X   VBGr�  G?�����X   CCr�  G?�7�7�X   NNr�  G?�{�{�X   MDr�  G?�����X   oovr�  G?�����X   JJr�  G?�*�*�X   NNPr�  G?���X   DTr�  G?�����X   NNSr�  G?���X   VBPr�  G?���X   VBDr�  G?�����X   NNPSr�  G?�����X   RBr�  G?�*�*�X   WDTr�  G?�����NG?�����X   WRBr�  G?���hMG?���X   TOr�  G?���uj)  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r   Rr  (X   NNr  G?�X   DTr  G?�X   JJr  G?�h�G?�X   PRP$r  G?�������X   VBNr  G?�UUUUUUX   TOr  G?�uX   JJr  hM�r	  h h(h
c__builtin__
__main__
hNN}r
  Ntr  Rr  �r  Rr  (X   ``r  G?��V��X   NNPr  G?��@�´HX   WPr  G?Ʒ*��
X   JJr  G?��$��X   CCr  G?�Ի~2z�X   WRBr  G?���{P�X   NNSr  G?�xm�|	X   DTr  G?��Ŗ�*�X   oovr  G?wxm�|	X   NNr  G?���{P�X   RBr  G?���{P�X   PRPr  G?�xm�|	X   INr  G?����vC�X   VBDr  G?�xm�|	X   CDr  G?�N�R5]X   ''r  G?�1	_��X   VBGr  G?��V��X   JJSr   G?wxm�|	X   VBr!  G?wxm�|	X   VBZr"  G?�N�R5]X   WDTr#  G?wxm�|	X   VBNr$  G?�N�R5]X   VBPr%  G?wxm�|	h�G?��V��X   TOr&  G?wxm�|	uj  j  �r'  h h(h
c__builtin__
__main__
hNN}r(  Ntr)  Rr*  �r+  Rr,  (X   NNPr-  G?�.:񍔄X   ''r.  G?���m��X   INr/  G?����|�YX   NNr0  G?����|�YX   VBZr1  G?�}�8��MX   RBr2  G?{��T�tX   TOr3  G?�}�8��Mh�G?�.:񍔄X   NNSr4  G?����>X   CCr5  G?���T�thMG?���T�tX   DTr6  G?r}�8��MX   RPr7  G?{��T�tX   POSr8  G?r}�8��MX   JJr9  G?{��T�tX   CDr:  G?r}�8��MX   ``r;  G?����+�2X   WRBr<  G?r}�8��MX   MDr=  G?r}�8��MX   VBDr>  G?r}�8��MuX   VBDr?  j�  �r@  h h(h
c__builtin__
__main__
hNN}rA  NtrB  RrC  �rD  RrE  (X   NNrF  G?�UUUUUUX   DTrG  G?�������X   NNPrH  G?ə�����X   VBGrI  G?�X   JJrJ  G?�X   CDrK  G?�X   VBNrL  G?�q�q�X   PRPrM  G?��l�lX   INrN  G?�q�q�X   NNSrO  G?��l�lX   VBrP  G?��l�lX   TOrQ  G?��l�lX   RBrR  G?��l�lX   oovrS  G?��l�lh�G?��l�lX   WPrT  G?��l�luX   VBDrU  j�  �rV  h h(h
c__builtin__
__main__
hNN}rW  NtrX  RrY  �rZ  Rr[  (X   WPr\  G?�/�A��4X   TOr]  G?ю���X   NNPr^  G?���!�xX   DTr_  G?���!�xX   NNr`  G?���!�xh�G?���!�xX   WRBra  G?���!�xX   VBGrb  G?�/�A��4X   PRPrc  G?�/�A��4X   INrd  G?���!�xX   VBNre  G?���ajzVX   MDrf  G?���!�xX   JJrg  G?���!�xX   PRP$rh  G?�/�A��4X   NNSri  G?�/�A��4X   RBrj  G?���!�xX   RPrk  G?���!�xX   oovrl  G?���!�xuj  j6  �rm  h h(h
c__builtin__
__main__
hNN}rn  Ntro  Rrp  �rq  Rrr  (X   VBDrs  G?��;�;h�G?͉؝�؞X   JJrt  G?�A�A�X   VBNru  G?�i�i�X   VBrv  G?��;�;X   RBrw  G?�A�A�X   NNrx  G?�i�i�X   INry  G?��;�;X   CCrz  G?�A�A�uj�  h��r{  h h(h
c__builtin__
__main__
hNN}r|  Ntr}  Rr~  �r  Rr�  NG?�      sj  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   CDr�  G?�`a�hX   NNSr�  G?�qj��&�X   DTr�  G?�Xo8�^X   NNPr�  G?���Ġh�G?����n-^X   VBGr�  G?���E�^X   INr�  G?��+���X   JJr�  G?���Ġ%X   PRP$r�  G?�D�d߳X   NNr�  G?�<ր(#�X   JJSr�  G?n�(�
�X   WPr�  G?�����X   PRPr�  G?�N�����X   RBr�  G?~�(�
�X   JJRr�  G?reЊѱ/X   TOr�  G?reЊѱ/X   VBPr�  G?`��O�[BX   VBDr�  G?yyw{�X   VBNr�  G?`��O�[BNG?gjO<P��X   VBZr�  G?Z£��^�X   WRBr�  G?n�(�
�X   oovr�  G?`��O�[BX   ``r�  G?Z£��^�X   WDTr�  G?d���X   NNPSr�  G?J£��^�X   CCr�  G?d���uX   INr�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   VBDr�  G?��<���\h�G?��R�7hMG?��:�YX   WRBr�  G?o��!ʩ�X   VBPr�  G?�~d��caX   WDTr�  G?�iu/W��X   VBZr�  G?�GQ��zX   INr�  G?�F�#�$PX   VBNr�  G?�H\mt$|X   TOr�  G?��s��X   POSr�  G?xR��;�iX   JJr�  G?���ǟX   ''r�  G?^��n<IQX   CCr�  G?����tg3X   MDr�  G?�iu/W��X   RBr�  G?��6aQ"X   NNSr�  G?�'C��v$X   CDr�  G?`��j��X   VBGr�  G?�u[��E�X   WPr�  G?��:�X   PRP$r�  G?@��j��X   NNr�  G?��_֐X   DTr�  G?m0	����X   NNPr�  G?v<�8��X   JJRr�  G?@��j��X   JJSr�  G?6<�8��X   PRPr�  G?V<�8��X   VBr�  G?o��!ʩ�X   oovr�  G?d�+�W�ZNG?F<�8��X   RBSr�  G?@��j��X   ``r�  G?F<�8��uX   JJr�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   NNr�  G?�[_u'X   WPr�  G?�[_u'X   INr�  G?�?�o^�X   DTr�  G?Æ�+c��X   JJr�  G?���/��X   VBr�  G?�[_u'X   VBNr�  G?���/��X   NNPr�  G?�$(F޼X   PRP$r�  G?���/��h�G?���/��X   TOr�  G?�[_u'X   VBGr�  G?�$(F޼X   NNSr�  G?�?�o^�X   RBr�  G?�$(F޼X   VBDr�  G?�[_u'X   VBPr�  G?�$(F޼X   RPr�  G?�[_u'X   PRPr�  G?��2��kX   WRBr�  G?�$(F޼hMG?�$(F޼uX   CDr�  j�
  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   WPr�  G?��O��X   RBr�  G?���`jc�X   VBr�  G?���C�X   CDr�  G?�7iH�X   DTr�  G?���`jc�X   NNPr�  G?��J@F�)h�G?��J@F�)X   JJr�  G?��J@F�)X   WRBr�  G?��J@F�)uj�
  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (h�G?�?
�yX   VBDr�  G?��+���X   INr�  G?��+���X   NNr�  G?��݄���X   JJr�  G?��b8l�]X   VBr�  G?���/9X   JJSr�  G?fJ�:��_X   NNSr�  G?����%��X   NNPr�  G?��b8l�hMG?����%��X   VBGr�  G?vJ�:��_X   VBZr�  G?��1Ί��X   MDr�  G?�J�:��_X   TOr�  G?fJ�:��_X   VBPr�  G?��8�8X   CDr�  G?��+���X   DTr   G?p���%��X   VBNr  G?fJ�:��_X   JJRr  G?fJ�:��_X   oovr  G?fJ�:��_X   RBr  G?fJ�:��_uX   ``r  j	  �r  h h(h
c__builtin__
__main__
hNN}r  Ntr  Rr	  �r
  Rr  (X   VBPr  G?ڪ�����X   VBZr  G?�������X   NNPSr  G?�      X   ''r  G?�      X   MDr  G?�UUUUUUX   VBDr  G?�      X   RBr  G?�UUUUUUX   WPr  G?�UUUUUUuj  j�  �r  h h(h
c__builtin__
__main__
hNN}r  Ntr  Rr  �r  Rr  (X   NNPr  G?�Ɉ+�WX   DTr  G?�W& �LAX   VBZr  G?�W& �LAX   VBNr  G?�W& �LX   INr  G?�W& �LX   CCr  G?�W& �LAX   JJr   G?�b
���X   VBDr!  G?�W& �LAX   RBr"  G?��;�6xX   NNr#  G?�Ɉ+�WX   NNSr$  G?�Ɉ+�WX   VBPr%  G?�Ɉ+�WX   PRPr&  G?�Ɉ+�Wuj�  j  �r'  h h(h
c__builtin__
__main__
hNN}r(  Ntr)  Rr*  �r+  Rr,  (X   NNPr-  G?�O1���X   NNSr.  G?�w�T�,4h�G?�ȿ�!'X   VBPr/  G?�ȿ�!'X   VBDr0  G?�BMZ>�cX   VBNr1  G?��V����X   oovr2  G?̋��j�hMG?�j����X   NNr3  G?��r/�X   CCr4  G?�ȿ�!&�X   INr5  G?�ȿ�!&�X   VBr6  G?�j����X   TOr7  G?�ȿ�!'X   POSr8  G?�j����X   ''r9  G?�j����X   DTr:  G?�ȿ�!'X   VBZr;  G?�w�T�,4X   RBr<  G?}w�T�,4X   CDr=  G?�ȿ�!'X   NNPSr>  G?}w�T�,4X   ``r?  G?}w�T�,4X   JJr@  G?}w�T�,4uX   VBNrA  j�  �rB  h h(h
c__builtin__
__main__
hNN}rC  NtrD  RrE  �rF  RrG  (h�G?��D��=�X   VBGrH  G?��D��=�X   JJrI  G?��D��=�X   PRPrJ  G?�
�B�P�X   INrK  G?�]�a�X   DTrL  G?�t�9GNX   NNPrM  G?���m�xX   NNSrN  G?����X   TOrO  G?���+@X   CDrP  G?����X   NNrQ  G?���m�xX   oovrR  G?����X   VBNrS  G?����X   RBrT  G?���+@X   WPrU  G?����X   CCrV  G?���+@X   VBDrW  G?���+@X   ``rX  G?���+@X   PRP$rY  G?���+@uX   VBrZ  h��r[  h h(h
c__builtin__
__main__
hNN}r\  Ntr]  Rr^  �r_  Rr`  (X   JJra  G?�������X   NNrb  G?��F#�X   NNSrc  G?��e��l�X   INrd  G?��w;���X   VBre  G?����X   CCrf  G?�������h�G?����X   TOrg  G?�
�B�P�X   RBrh  G?����X   WPri  G?�
�B�P�X   VBNrj  G?�
�B�P�uh�ja  �rk  h h(h
c__builtin__
__main__
hNN}rl  Ntrm  Rrn  �ro  Rrp  (X   NNrq  G?�UUUUUUX   NNPrr  G?�X   NNSrs  G?�g�g�h�G?��p�pX   CCrt  G?�X   INru  G?��?��?�X   WRBrv  G?��p�phMG?��p�pX   TOrw  G?��f�fX   JJrx  G?�X   oovry  G?��p�puX   VBDrz  j�  �r{  h h(h
c__builtin__
__main__
hNN}r|  Ntr}  Rr~  �r  Rr�  (X   NNPr�  G?����X   INr�  G?�De�JBX   ``r�  G?t�C��,LX   PRP$r�  G?�T��7^X   DTr�  G?�JBqW�^X   WRBr�  G?De�JBqX   RBr�  G?�T��7^h�G?�=;G ��X   JJr�  G?��C��,LX   WPr�  G?��]&n��hMG?��C��,LX   VBGr�  G?�%����X   NNSr�  G?�����i�X   NNr�  G?�=;G ��X   WDTr�  G?De�JBqX   CCr�  G?t�C��,LX   JJSr�  G?��C��,LX   CDr�  G?��C��,LX   TOr�  G?�sL6���uj�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   INr�  G?��8�8X   NNPr�  G?�ѭѭh�G?��_�_X   CCr�  G?�A�A�X   POSr�  G?�)r�)r�X   NNSr�  G?�a�a�X   NNr�  G?�A�A�X   RBr�  G?��8�8X   VBZr�  G?��8�8X   VBPr�  G?��8�8uj  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   WRBr�  G?�Q���4X   VBNr�  G?�e���X   PRPr�  G?�`�vO��X   INr�  G?��p0��X   RBr�  G?���򽴇X   NNr�  G?�[����X   DTr�  G?�`�vO��X   WPr�  G?�[����X   NNPr�  G?�e���h�G?�zc���X   TOr�  G?�Q���4X   PRP$r�  G?�p0���X   WDTr�  G?�zc���X   JJr�  G?�V�wT�DX   NNSr�  G?����X   RPr�  G?�zc���X   oovr�  G?�Q���4X   VBGr�  G?�Q���4uh\j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   DTr�  G?��"Gy��X   INr�  G?�>�@�c�X   VBGr�  G?�r�LV��X   PRP$r�  G?�,}r���X   TOr�  G?��6u.oYh�G?�q�q�X   NNSr�  G?���X   NNPr�  G?���˺�X   RPr�  G?�]פ��3X   NNr�  G?�,}r���hMG?c�WG<X   RBr�  G?�c�WG<X   VBNr�  G?�k�i�F�X   PRPr�  G?�,}r���X   JJr�  G?����7X   oovr�  G?gV��umX   VBr�  G?{:�7�^TX   WRBr�  G?�V��umX   CCr�  G?oc�WG<X   WPr�  G?oc�WG<X   MDr�  G?gV��umX   ``r�  G?�V��umX   RBSr�  G?_c�WG<X   VBZr�  G?oc�WG<X   CDr�  G?sr�LV��X   VBDr�  G?_c�WG<X   JJRr�  G?_c�WG<X   WDTr�  G?_c�WG<uX   WRBr�  h?�r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   VBDr�  G?��x�g�jX   oovr�  G?���؍wX   INr�  G?���؍wnX   RPr�  G?j��؍wh�G?�Ú�	�9X   VBZr�  G?ǫ��@4X   PRPr�  G?qiH�;�X   VBNr�  G?��q��jX   JJRr�  G?�K	?�X   RBr�  G?�ey�WTX   VBPr�  G?�#����X   MDr�  G?�|%��X   CDr�  G?uÚ�	�9X   TOr�  G?j��؍wX   JJr�  G?z��؍wX   DTr�  G?�iH�;�X   VBGr�  G?qiH�;�X   NNr�  G?qiH�;�uX   NNr�  j  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   INr�  G?�lߡ���X   DTr�  G?˞�	\��X   NNr�  G?����Z&X   RPr�  G?��F�`�X   NNPr�  G?��+��fX   JJSr�  G?y�$�U�X   RBr�  G?�I8�a�X   VBNr�  G?�I8�a�h�G?�I8�a�X   JJr�  G?���%��8X   NNSr   G?�&ɲl�'X   TOr  G?��8����X   JJRr  G?�0�{Q��X   CDr  G?�ft�8�X   RBSr  G?���,�E�X   WPr  G?��ռ��X   PRPr  G?���S1|�X   PRP$r  G?���|X   WDTr  G?eft�8�X   VBGr	  G?�B���̤X   VBr
  G?sB���̤X   NNPSr  G?m�ռ��X   CCr  G?Y�$�U�X   VBZr  G?{��S1|�X   VBDr  G?uft�8�NG?Y�$�U�X   ``r  G?Q�F�`�hMG?Q�F�`�X   WRBr  G?sB���̤X   oovr  G?eft�8�X   MDr  G?Q�F�`�uX   NNr  je  �r  h h(h
c__builtin__
__main__
hNN}r  Ntr  Rr  �r  Rr  (X   VBr  G?��GF��X   DTr  G?�'��nX   NNr  G?��*�`X   RBr  G?���ϰ��X   NNSr  G?�����YKX   NNPr  G?�����YKX   CDr   G?��:5u�X   PRPr!  G?��0�@X�X   VBGr"  G?c�*�`hMG?YW��Z��h�G?s�*�`X   INr#  G?c�*�`X   PRP$r$  G?YW��Z��X   JJr%  G?s�*�`X   ``r&  G?iW��Z��uj  j`  �r'  h h(h
c__builtin__
__main__
hNN}r(  Ntr)  Rr*  �r+  Rr,  (X   TOr-  G?�������X   INr.  G?�������X   DTr/  G?ə�����X   RBr0  G?�333333X   VBNr1  G?�������X   NNPr2  G?�      X   JJr3  G?�������X   WDTr4  G?�������X   ``r5  G?�������X   WPr6  G?�������X   PRP$r7  G?�������X   NNSr8  G?�������uj�  ja  �r9  h h(h
c__builtin__
__main__
hNN}r:  Ntr;  Rr<  �r=  Rr>  (X   NNPr?  G?Ê��!!�X   INr@  G?���B� �X   NNrA  G?� �R�+�X   NNSrB  G?��Dmϕ�X   VBNrC  G?�:k��@�X   DTrD  G?ӭ<s8d�X   CDrE  G?�dX,[kh�G?�Ob�U�X   VBGrF  G?�<P���'X   PRPrG  G?�W��Z��X   JJrH  G?��H7-�X   VBrI  G?�Ob�U�X   WPrJ  G?�dX,[kX   PRP$rK  G?��p��K�X   oovrL  G?nJ�ZVHX   WRBrM  G?�dX,[k>hMG?aOb�U�X   RBrN  G?w�&���X   WDTrO  G?syNM��X   ``rP  G?w�&���X   TOrQ  G?~J�ZVHX   JJSrR  G?e�:���XX   NNPSrS  G?QOb�U�X   VBDrT  G?aOb�U�X   CCrU  G?Y�r �X   JJRrV  G?e�:���XX   MDrW  G?QOb�U�uhMj*  �rX  h h(h
c__builtin__
__main__
hNN}rY  NtrZ  Rr[  �r\  Rr]  (hMG?���|h�G?�q�q�X   INr^  G?�l�&ɲmX   TOr_  G?��֠R�[X   NNSr`  G?��֠R�[X   CCra  G?��֠R�[X   NNrb  G?���Hgo1X   NNPrc  G?��֠R�[X   RBrd  G?��֠R�[uj*  hM�re  h h(h
c__builtin__
__main__
hNN}rf  Ntrg  Rrh  �ri  Rrj  (X   INrk  G?���s���X   VBDrl  G?����X   WPrm  G?ш�b1�X   WRBrn  G?���s���X   CDro  G?�
�B�P�X   RBrp  G?��F#��X   VBNrq  G?�
�B�P�X   CCrr  G?��F#��X   NNSrs  G?�
�B�P�X   WDTrt  G?���b1�X   DTru  G?��F#��X   JJrv  G?����X   PRPrw  G?����X   NNrx  G?����X   VBGry  G?���b1�X   NNPrz  G?����X   VBZr{  G?����X   TOr|  G?�
�B�P�X   MDr}  G?����uj}
  j.  �r~  h h(h
c__builtin__
__main__
hNN}r  Ntr�  Rr�  �r�  Rr�  (X   VBDr�  G?�,I���X   NNPr�  G?�������h�G?�����:XX   NNr�  G?�N�$�`X   CCr�  G?��u�
�^X   RBr�  G?��u�
�^X   CDr�  G?�0ѐX   NNPSr�  G?�����:XX   VBZr�  G?�����:XX   MDr�  G?�0ѐX   VBPr�  G?��_A}�X   JJr�  G?�����:XX   POSr�  G?�0ѐhMG?s0ѐX   TOr�  G?|����:XX   INr�  G?��_A}�X   NNSr�  G?��u�
�^X   VBNr�  G?|����:XX   VBr�  G?s0ѐuX   NNr�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   VBDr�  G?��vr�X   VBPr�  G?�&5~��X   VBZr�  G?��g*�LX   INr�  G?�H���\X   MDr�  G?���[��X   NNr�  G?���@�X   TOr�  G?��vr�zX   RBr�  G?���@�X   JJSr�  G?~�1��gh�G?�1��g*X   NNPr�  G?��1��gX   DTr�  G?��vr�zhMG?���@�X   VBr�  G?~�1��gX   JJr�  G?���@�X   VBNr�  G?~�1��gX   ''r�  G?~�1��gX   NNSr�  G?��1��gX   VBGr�  G?~�1��gX   ``r�  G?���@�uX   INr�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (h�G?���g*X   NNSr�  G?��[���X   TOr�  G?�H���\X   INr�  G?�r�zDưX   JJr�  G?��vr�zX   VBNr�  G?��vr�zX   NNr�  G?ĉ�_��9X   VBZr�  G?��vr�X   CCr�  G?���@�X   CDr�  G?���@�X   VBDr�  G?��1��gX   RBr�  G?��1��gX   NNPr�  G?��1��gX   DTr�  G?���@�X   POSr�  G?~�1��gX   WPr�  G?~�1��gX   RPr�  G?���@�X   JJRr�  G?���@�uX   RBr�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   INr�  G?��y�u�X   VBDr�  G?�.)��GXX   DTr�  G?�.)��GXX   JJr�  G?�d���mX   VBNr�  G?�.)��GXX   NNr�  G?��ͣ�X   VBr�  G?�`�K�}�X   RBr�  G?��ͣ��X   CDr�  G?�.)��GXX   NNSr�  G?��qO��;X   CCr�  G?��qO��;hMG?��qO��;X   VBZr�  G?�.)��GXX   JJRr�  G?��qO��;X   WPr�  G?��qO��;X   NNPSr�  G?��qO��;uX   JJSr�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   INr�  G?�󯢬eh�G?�Mū�0�X   NNr�  G?�3�* hX   VBDr�  G?�qj��&�X   VBPr�  G?��Ly��VX   RBr�  G?�쎕3�X   ''r�  G?�Ly��hMG?��Ly��X   WRBr�  G?��>ݦ��X   VBGr�  G?��>ݦ��X   VBNr�  G?��Ly��X   RPr�  G?t�>ݦ��X   WDTr�  G?��>ݦ��X   VBr�  G?t�>ݦ��X   TOr�  G?���T�X   WPr�  G?t�>ݦ��X   CCr�  G?�쎕3�X   VBZr�  G?t�>ݦ��X   NNSr�  G?��>ݦ��X   DTr�  G?t�>ݦ��X   NNPr�  G?t�>ݦ��X   JJr�  G?��>ݦ��X   MDr�  G?t�>ݦ��uX   CDr�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   VBDr�  G?�����/hX   INr   G?�H�����X   VBNr  G?��<�X~X   NNr  G?�H�����X   WRBr  G?�H�����X   TOr  G?�����/hX   RBr  G?�����/hX   NNSr  G?�H�����X   DTr  G?�����/hX   VBZr  G?�H�����X   JJr	  G?���<�XX   WPr
  G?�H�����X   PRPr  G?�H�����X   NNPr  G?���<�Xh�G?�����/hX   JJRr  G?�H�����X   oovr  G?�H�����X   RBSr  G?�H�����uj�  j�  �r  h h(h
c__builtin__
__main__
hNN}r  Ntr  Rr  �r  Rr  (X   NNPr  G?Ӆ���BX   INr  G?��`����X   DTr  G?�-�JX   VBNr  G?� 3����X   PRPr  G?�R�+x�X   NNSr  G?���N�X   RPr  G?�R�+x�X   TOr  G?�&�9�V�X   NNr  G?���N�X   JJr  G?���N�X   RBr   G?���N�X   oovr!  G?y��N�X   VBr"  G?�R�+x�X   CCr#  G?y��N�X   RBSr$  G?y��N�X   JJRr%  G?y��N�X   VBGr&  G?y��N�X   NNPSr'  G?y��N�X   PRP$r(  G?�R�+x�uh�jb  �r)  h h(h
c__builtin__
__main__
hNN}r*  Ntr+  Rr,  �r-  Rr.  (X   INr/  G?�ƥ/�X   RPr0  G?�/�a�jX   TOr1  G?�a�jQ"�X   PRP$r2  G?��H�@Y�X   WPr3  G?��0�5)X   JJr4  G?��y�u�X   NNSr5  G?�d���mX   DTr6  G?��=�J$X   NNPr7  G?�a�jQ"�X   VBGr8  G?�a�jQ"�X   oovr9  G?{�g��k�X   VBr:  G?p�qO��;X   RBr;  G?��ͣ��X   WRBr<  G?������h�G?�d���mX   NNr=  G?�H�@Y��X   VBNr>  G?�.)��GXX   JJSr?  G?p�qO��;X   VBPr@  G?fa�jQ"�X   CDrA  G?{�g��k�X   CCrB  G?va�jQ"�X   JJRrC  G?������X   PRPrD  G?�a�jQ"�X   VBZrE  G?fa�jQ"�X   WDTrF  G?p�qO��;hMG?fa�jQ"�X   VBDrG  G?fa�jQ"�X   ``rH  G?p�qO��;NG?fa�jQ"�uX   WPrI  j�  �rJ  h h(h
c__builtin__
__main__
hNN}rK  NtrL  RrM  �rN  RrO  (X   JJSrP  G?}e�B$�X   DTrQ  G?�]E�t]X   NNPrR  G?Ù,cX   VBGrS  G?�?���PX   CDrT  G?�%���owX   INrU  G?��,cX   PRP$rV  G?�,c7X   JJrW  G?�����'2X   NNSrX  G?�����3rX   NNrY  G?���ǧ�X   VBNrZ  G?}e�B$�X   TOr[  G?s�,cX   PRPr\  G?�e�B$�X   VBZr]  G?s�,cX   WDTr^  G?s�,cX   RBr_  G?}e�B$�X   VBDr`  G?s�,cX   JJRra  G?s�,cX   NNPSrb  G?}e�B$�h�G?s�,cuX   WPrc  j
  �rd  h h(h
c__builtin__
__main__
hNN}re  Ntrf  Rrg  �rh  Rri  (X   VBDrj  G?�t�j �X   VBZrk  G?�'�᭲�X   RBrl  G?�ʸ�%�nX   VBNrm  G?��G�(�h�G?�d�
eX   JJrn  G?�)&�6%X   NNSro  G?{��	���X   INrp  G?�S�����X   VBPrq  G?�����r�X   MDrr  G?�ʸ�%�nX   VBGrs  G?k��	���X   VBrt  G?k��	���X   CCru  G?k��	���NG?k��	���hMG?�A�HV�X   NNPrv  G?k��	���X   WRBrw  G?k��	���X   TOrx  G?k��	���X   NNry  G?k��	���uX   RBSrz  jW  �r{  h h(h
c__builtin__
__main__
hNN}r|  Ntr}  Rr~  �r  Rr�  (X   INr�  G?�$�I$�IX   RBr�  G?�m��m��X   VBGr�  G?�I$�I$�X   VBPr�  G?�$�I$�Ih�G?ВI$�I%X   WRBr�  G?�I$�I$�X   VBDr�  G?�I$�I$�X   VBr�  G?�I$�I$�X   CCr�  G?�m��m��X   VBNr�  G?�      X   TOr�  G?�I$�I$�X   POSr�  G?�I$�I$�X   NNSr�  G?�I$�I$�X   DTr�  G?�I$�I$�X   NNr�  G?�I$�I$�uX   RBSr�  jX  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   NNSr�  G?��8�9X   NNPr�  G?��q�rX   VBZr�  G?�q�q�X   VBr�  G?�q�q�X   VBPr�  G?�q�q�X   VBDr�  G?�q�q�X   JJr�  G?�q�q�X   NNr�  G?�UUUUUUh�G?�q�q�X   NNPSr�  G?�UUUUUUX   INr�  G?�q�q�uX   RBSr�  jY  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   CDr�  G?�򆼡�(X   INr�  G?ܡ�(k�h�G?�Pה5�X   TOr�  G?�ה5�yX   NNSr�  G?��5�yCX   VBNr�  G?�5�yC^X   NNr�  G?�5�yC^X   CCr�  G?�򆼡�(X   VBGr�  G?�򆼡�(X   VBPr�  G?�򆼡�(X   RBr�  G?�򆼡�(uX   VBZr�  j   �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   CDr�  G?��Aq�X   WPr�  G?��g��&X   DTr�  G?�i9NF�X   NNSr�  G?�WBЅX   NNPr�  G?�pG��h�G?���屹lX   PRP$r�  G?��}�pX   VBGr�  G?�򆼡�(X   oovr�  G?��}�pX   WDTr�  G?���+�
�X   WRBr�  G?~����X   JJr�  G?�3T�5X   INr�  G?��"H�X   VBDr�  G?n����X   NNr�  G?�gLY�uX   VBPr�  G?^����X   JJSr�  G?t�"H�X   PRPr�  G?��j���X   TOr�  G?w�Aq�X   ``r�  G?|;�ðX   CCr�  G?q�}�pX   VBZr�  G?i�j���X   RBr�  G?|;�ðX   ''r�  G?T�"H�X   VBNr�  G?t�"H�X   VBr�  G?T�"H�X   JJRr�  G?t�"H�NG?T�"H�X   NNPSr�  G?^����hMG?^����uX   CCr�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   JJr�  G?�      X   NNr�  G?�      X   NNSr�  G?�      X   WPr�  G?�      X   VBNr�  G?�      X   NNPr�  G?�      uj�  hÆr�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   NNr�  G?�Me5��SX   DTr�  G?��_A}�X   TOr�  G?��_A}�X   NNSr�  G?��/���X   JJr�  G?Ŕ�SYMeX   JJRr�  G?��_A}�X   POSr�  G?��_A}�h�G?��_A}�X   VBNr�  G?��Gq�wuX   VBDr�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   INr�  G?�lB:�I�X   WRBr�  G?qw�քX   VBPr�  G?��1��gX   VBGr�  G?�3O%���X   VBDr�  G?��{\?QUX   TOr�  G?��9�eX?X   RBr�  G?��ԃ��X   VBNr�  G?�x���C�X   CDr�  G?m�ԃ��X   VBr�  G?�xDi��X   MDr�  G?gJv�Ȱh�G?��A���X   CCr   G?�b@h�<�X   NNr  G?���@:9"X   oovr  G?wJv�ȰX   JJr  G?��A���X   DTr  G?�w�քX   NNSr  G?wJv�ȰhMG?}�ԃ��X   POSr  G?wJv�ȰX   WPr  G?t`���ϚX   WDTr  G?�����QX   VBZr	  G?t`���ϚX   PRPr
  G?aw�քX   NNPr  G?m�ԃ��X   JJSr  G?WJv�ȰNG?WJv�ȰX   JJRr  G?gJv�ȰX   RPr  G?WJv�ȰX   ''r  G?aw�քujv  j�  �r  h h(h
c__builtin__
__main__
hNN}r  Ntr  Rr  �r  Rr  (X   NNPr  G?�+n6���X   VBGr  G?��O8�.X   PRPr  G?��� o��X   CDr  G?��0��<X   PRP$r  G?��`v���X   DTr  G?�&�^HX   INr  G?��b�L�X   NNr  G?�>��T�X   WPr  G?�Uv��X   WDTr  G?�u�'�j�X   WRBr   G?��� o��h�G?��`v���X   TOr!  G?k�i�'�X   JJr"  G?���l�V�X   VBDr#  G?[�i�'�X   NNSr$  G?��1�t�X   JJRr%  G?t�b�L�X   VBZr&  G?d�b�L�X   oovr'  G?[�i�'�X   NNPSr(  G?[�i�'�X   JJSr)  G?d�b�L�X   CCr*  G?[�i�'�X   VBr+  G?[�i�'�X   VBNr,  G?[�i�'�X   RBr-  G?d�b�L�uX   TOr.  j�  �r/  h h(h
c__builtin__
__main__
hNN}r0  Ntr1  Rr2  �r3  Rr4  (X   INr5  G?�����/hX   NNSr6  G?Ǵ%�	{BX   JJr7  G?�����/hX   CCr8  G?�����/hX   NNr9  G?�����/hX   RBr:  G?�����/hX   DTr;  G?�����/huX   NNr<  j  �r=  h h(h
c__builtin__
__main__
hNN}r>  Ntr?  Rr@  �rA  RrB  (X   NNSrC  G?�X   NNrD  G?ᱱ����h�G?�X   JJrE  G?�X   JJSrF  G?�X   RBrG  G?�X   INrH  G?�X   CDrI  G?�X   TOrJ  G?�X   ``rK  G?�ujC  j�  �rL  h h(h
c__builtin__
__main__
hNN}rM  NtrN  RrO  �rP  RrQ  (h�G?�T:�)X   VBrR  G?�W�p\C�X   WPrS  G?����X   PRP$rT  G?��B��cX   NNSrU  G?��R�g��X   INrV  G?y)É�cX   NNPrW  G?���mX   DTrX  G?Ğ��PcX   NNrY  G?�^%8q<X   VBGrZ  G?���W��PX   JJr[  G?�[d ��X   CCr\  G?`Ƃ[�T�X   WRBr]  G?s�B��cX   WDTr^  G?�Ƃ[�T�X   CDr_  G?`Ƃ[�T�X   ``r`  G?s�B��cX   RBra  G?~�DS-��X   oovrb  G?f^%8q<X   JJSrc  G?`Ƃ[�T�X   JJRrd  G?V^%8q<X   VBNre  G?V^%8q<X   PRPrf  G?v^%8q<hMG?V^%8q<X   NNPSrg  G?V^%8q<uX   NNrh  j�  �ri  h h(h
c__builtin__
__main__
hNN}rj  Ntrk  Rrl  �rm  Rrn  (h�G?�)����UX   VBro  G?`$6Qz7X   DTrp  G?�':�Df�X   NNPrq  G?�!1ʰX   INrr  G?��S};��X   VBNrs  G?Ȥ�s,�%X   TOrt  G?�%���N�X   NNru  G?�.�)=��X   PRP$rv  G?���X	X   WPrw  G?x$6Qz7SX   JJrx  G?�%���N�X   RPry  G?�':�Df�X   RBrz  G?�$6Qz7SX   VBGr{  G?�-C���X   PRPr|  G?t-C���X   NNSr}  G?�(��~X   WRBr~  G?�-C���X   JJRr  G?�(��~hMG?`$6Qz7X   oovr�  G?p$6Qz7X   JJSr�  G?h$6Qz7SX   WDTr�  G?`$6Qz7NG?`$6Qz7X   CCr�  G?`$6Qz7X   VBDr�  G?h$6Qz7SX   CDr�  G?h$6Qz7SX   ``r�  G?`$6Qz7uX   VBr�  h��r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   INr�  G?�E�t]Fh�G?�E�t]X   TOr�  G?���|hMG?�E�t]FX   VBr�  G?�6M�d�6X   JJr�  G?����>�X   VBPr�  G?�d�6M�eX   CDr�  G?�d�6M�eX   CCr�  G?�&ɲl�'X   VBNr�  G?��>���X   NNPr�  G?��|X   RBr�  G?�>���>X   DTr�  G?�l�&ɲmX   ''r�  G?o��|X   WPr�  G?wE�t]FX   NNr�  G?�d�6M�eX   JJRr�  G?�&ɲl�'X   oovr�  G?�d�6M�eX   PRPr�  G?wE�t]FX   NNSr�  G?wE�t]FX   VBGr�  G?�E�t]FX   WRBr�  G?o��|X   ``r�  G?o��|uX   VBr�  j   �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   INr�  G?��j�(X   PRPr�  G?����MX   VBZr�  G?�����;�X   NNr�  G?̛�ueh�G?�\�o��X   TOr�  G?��}���+X   CDr�  G?��R_�9X   RBr�  G?����;�X   NNPr�  G?����;�X   JJr�  G?��e�\�pX   NNSr�  G?��R_�9X   DTr�  G?����;�X   VBDr�  G?����;�X   VBr�  G?��"���NG?w�"���X   MDr�  G?o����;�X   CCr�  G?o����;�X   VBNr�  G?o����;�hMG?w�"���uX   NNSr�  j=  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (h�G?�a�a�X   NNPr�  G?�a�a�X   INr�  G?�UUUUUUX   VBGr�  G?�UUUUUUX   VBr�  G?�a�a�X   PRPr�  G?�m��m��X   NNr�  G?�a�a�X   DTr�  G?�0�0�X   RBr�  G?�a�a�X   VBNr�  G?��<��<�X   NNSr�  G?�I$�I$�X   WDTr�  G?�a�a�X   VBZr�  G?�a�a�X   JJr�  G?�m��m��X   WPr�  G?�I$�I$�X   VBDr�  G?�I$�I$�X   CDr�  G?�a�a�NG?�a�a�X   NNPSr�  G?�a�a�X   TOr�  G?�I$�I$�X   VBPr�  G?�a�a�X   oovr�  G?�I$�I$�uj�  h��r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (NG?��5F�X   ``r�  G?l�\��y X   NNr�  G?l�\��y uX   VBDr�  h]�r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   VBNr�  G?r��+@X   NNSr�  G?�I��i4�X   JJr�  G?��Ƹ��,X   INr�  G?ՠ%h	ZX   NNr�  G?�a�Avh�G?��D��=�X   NNPr�  G?�]�a�X   CCr�  G?�]�a�X   RBr�  G?r��+@X   WPr�  G?r��+@X   TOr�  G?���+@X   POSr�  G?|���X   CDr�  G?���b1�hMG?�]�a�X   DTr�  G?�a�AvX   NNPSr�  G?r��+@X   ''r�  G?r��+@X   JJRr�  G?r��+@uh]j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (h�G?�SjmM��X   INr�  G?�jmM��7X   TOr�  G?�"�P�BX   VBNr�  G?��\�pX   WPr�  G?��\�pX   VBDr�  G?��\�pX   NNr�  G?�B(E�X   WDTr   G?��\�pX   NNSr  G?��\�pX   JJr  G?��\�puX   PRP$r  j�  �r  h h(h
c__builtin__
__main__
hNN}r  Ntr  Rr  �r  Rr	  (X   NNr
  G?�UUUUUUX   NNSr  G?�UUUUUUujY
  j�  �r  h h(h
c__builtin__
__main__
hNN}r  Ntr  Rr  �r  Rr  (X   INr  G?�f�NK�wX   JJr  G?����R#X   NNPr  G?�T�S��X   VBNr  G?��c�DQ^X   DTr  G?�IN�?�OX   PRPr  G?��c�DQX   TOr  G?�l;�8X   NNSr  G?��O�tKX   PRP$r  G?��Yϣ��X   RPr  G?��c�DQ^X   WPr  G?�J׳=X   NNr  G?�	��n�gX   NNPSr  G?rl;�8h�G?��c�DQ^X   WRBr  G?��c�DQ^X   CCr   G?�l;�8X   VBGr!  G?��6�r_�X   JJSr"  G?~�c�DQ^X   oovr#  G?rl;�8X   RBr$  G?�J׳=X   WDTr%  G?rl;�8X   CDr&  G?~�c�DQ^X   JJRr'  G?x�O�tKX   VBr(  G?rl;�8X   ``r)  G?��O�tKX   VBDr*  G?h�O�tKujN	  j�  �r+  h h(h
c__builtin__
__main__
hNN}r,  Ntr-  Rr.  �r/  Rr0  (X   JJr1  G?�#Or�4�X   NNr2  G?��i�XGX   NNSr3  G?ǹa{�X   VBGr4  G?���a|X   NNPr5  G?���a{�X   VBNr6  G?�{���aX   WPr7  G?���a{�X   JJSr8  G?�{���aX   ``r9  G?���a{�uX   NNr:  j  �r;  h h(h
c__builtin__
__main__
hNN}r<  Ntr=  Rr>  �r?  Rr@  (X   VBNrA  G?�F�]�h�G?{������X   NNPrB  G?�߭T�B�X   WRBrC  G?qț?lX   PRPrD  G?����L=�X   RBrE  G?�Pά�X�X   WPrF  G?�̱�+X   DTrG  G?�%}b�@X   VBDrH  G?h+��q~X   ``rI  G?t/���6_X   INrJ  G?��c!�klX   VBrK  G?���u�~�X   VBGrL  G?�Q� ��X   JJrM  G?�wB%٫JX   JJRrN  G?w�1b�X   TOrO  G?��ң�[X   PRP$rP  G?qM�!�
	X   NNrQ  G?���nɂX   oovrR  G?x�A���EX   CDrS  G?�ԏ��X   VBZrT  G?`Wy���AX   RBSrU  G?w�1b�X   RPrV  G?rC�\g�X   WDTrW  G?X�A���EX   NNSrX  G?�ey���8hMG?S9��)'�X   CCrY  G?G�1b�X   VBPrZ  G?S9��)'�X   JJSr[  G?i�X2w�NG?>��XA��X   NNPSr\  G?>��XA��X   POSr]  G?7�1b�X   ''r^  G?.��XA��uj  jA  �r_  h h(h
c__builtin__
__main__
hNN}r`  Ntra  Rrb  �rc  Rrd  (X   WPre  G?�o;�%�bX   INrf  G?�J3qA-X   WDTrg  G?^*H�,	(X   NNPrh  G?���]R��X   VBNri  G?��ܕ5�RX   JJrj  G?��[M��qX   TOrk  G?�0�J3qAX   NNrl  G?�P��HsFX   DTrm  G?���h�'X   VBGrn  G?�������h�G?�.FK��X   RBro  G?� ���X   RPrp  G?�ơ�U`�hMG?w��}�+�X   JJRrq  G?n*H�,	(X   WRBrr  G?���h�'X   NNSrs  G?�)���QX   PRP$rt  G?^*H�,	(X   oovru  G?n*H�,	(X   CCrv  G?v�����X   CDrw  G?e������X   JJSrx  G?U������X   RBSry  G?a<��bN`X   PRPrz  G?e������X   VBDr{  G?U������X   VBZr|  G?U������X   VBr}  G?^*H�,	(NG?A<��bN`X   ''r~  G?I���u�X   MDr  G?A<��bN`X   ``r�  G?Y���u�uX   RBr�  h��r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (NG?�4V�YX   ''r�  G?k�y�3X   ``r�  G?[�y�3X   NNPr�  G?[�y�3X   NNSr�  G?[�y�3X   CCr�  G?dB��}&�uX   TOr�  j   �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   NNr�  G?۠�lz�X   JJr�  G?ƾ'ڹ�X   VBZr�  G?O�$�K�0X   CDr�  G?�UEu��X   NNSr�  G?������[X   NNPr�  G?�L�V5�X   VBNr�  G?�P�MբX   VBGr�  G?{�@
�a�X   WPr�  G?bd*��AX   JJSr�  G?e�2�uX   DTr�  G?bd*��AX   JJRr�  G?vUEu��X   NNPSr�  G?���Tg]X   RBr�  G?rd*��AX   ``r�  G?bd*��AX   INr�  G?���
�kh�G?o�$�K�0X   VBDr�  G?E�2�uX   oovr�  G?_�$�K�0hMG?U�2�uX   RBSr�  G?E�2�uX   WDTr�  G?E�2�uX   VBr�  G?E�2�uX   WRBr�  G?E�2�uuX   INr�  jM  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   NNr�  G?�m`�K�X   NNPr�  G?��ͣ��X   VBZr�  G?�.)��GXX   JJr�  G?�GX!��X   DTr�  G?��ͣ�X   CDr�  G?��ͣ��X   MDr�  G?��qO��;X   RBr�  G?��ͣ��X   VBDr�  G?��d���X   INr�  G?��qO��;X   NNSr�  G?��ͣ�X   VBPr�  G?��qO��;X   CCr�  G?�.)��GXX   oovr�  G?�.)��GXh�G?��qO��;X   VBGr�  G?��qO��;NG?��qO��;ujM  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   VBDr�  G?ə�����X   NNPr�  G?�W:��tX   INr�  G?���j1M�h�G?�-��-��hMG?�W:��tX   oovr�  G?��So��X   VBZr�  G?�����/hX   CCr�  G?�W:��tX   NNr�  G?�W:��X   CDr�  G?�W:��tX   MDr�  G?��l�lX   VBPr�  G?�����/hX   TOr�  G?�����/hX   ''r�  G?�����/hX   VBGr�  G?��l�lX   RBr�  G?��l�lX   NNSr�  G?�����/hX   VBNr�  G?�W:��tX   WDTr�  G?~W:��tX   PRPr�  G?~W:��tX   DTr�  G?�W:��tX   JJr�  G?~W:��tuj  jo  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (h�G?�I�1@ �X   NNr�  G?�V��"X   INr�  G?��`r��GX   DTr�  G?�6ay�QX   TOr�  G?���c�X   NNPr�  G?����&zX   PRPr�  G?������8X   RBr�  G?�xP5[X   RPr�  G?������8X   VBNr�  G?�ο�*��X   VBr�  G?�xP5[X   WPr�  G?�j��y�X   VBGr�  G?��j��yX   PRP$r�  G?��j��yX   JJr�  G?��I\ۓX   CDr�  G?x�j��yX   WDTr�  G?x�j��yX   NNSr�  G?��c�W�X   JJSr�  G?x�j��yX   WRBr�  G?pj��y�X   VBZr�  G?pj��y�X   POSr�  G?pj��y�X   CCr�  G?pj��y�X   oovr�  G?pj��y�X   ''r�  G?pj��y�X   ``r�  G?x�j��yuX   POSr�  jR  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   DTr   G?�������X   JJr  G?�X   NNr  G?�������X   VBPr  G?�X   NNPr  G?ׇ�����X   INr  G?�X   MDr  G?�X   oovr  G?�X   VBDr  G?�X   NNSr	  G?�X   VBGr
  G?�X   WRBr  G?�X   CDr  G?�uNh(�r  h h(h
c__builtin__
__main__
hNN}r  Ntr  Rr  �r  Rr  (X   INr  G?�X��Ƈ�X   NNr  G?�
r�S��X   CCr  G?�X��ƈX   JJr  G?���/9X   VBZr  G?���/9X   NNPr  G?�X��ƈX   NNSr  G?ǂ����hMG?���/9X   VBDr  G?���/9X   MDr  G?���/9uX   POSr  jS  �r  h h(h
c__builtin__
__main__
hNN}r  Ntr  Rr   �r!  Rr"  (X   JJr#  G?�}}}}}}X   NNPr$  G?�X   NNSr%  G?�uX   NNPr&  h��r'  h h(h
c__builtin__
__main__
hNN}r(  Ntr)  Rr*  �r+  Rr,  (X   NNr-  G?�Ƹ-��X   INr.  G?�Q�����X   TOr/  G?��W> �X   VBDr0  G?��Q�<]h�G?����q�X   NNSr1  G?�ː��X   JJr2  G?���8f9HX   RBr3  G?�3��yX   NNPr4  G?�M�����X   VBPr5  G?�&Uz���X   NNPSr6  G?l3��yX   PRPr7  G?\3��yX   VBGr8  G?u&Uz���X   VBZr9  G?u&Uz���X   CCr:  G?�o�٪�X   VBNr;  G?��8f9HhMG?u&Uz���X   ``r<  G?\3��yX   ''r=  G?\3��yX   RPr>  G?\3��yX   VBr?  G?e&Uz���X   CDr@  G?u&Uz���X   WDTrA  G?\3��yX   JJRrB  G?\3��yX   WRBrC  G?\3��yuj	  h��rD  h h(h
c__builtin__
__main__
hNN}rE  NtrF  RrG  �rH  RrI  NG?�      sX   oovrJ  j�  �rK  h h(h
c__builtin__
__main__
hNN}rL  NtrM  RrN  �rO  RrP  (X   PRP$rQ  G?��L�x��X   NNPrR  G?��L�x��X   RPrS  G?���a{�X   RBrT  G?�{���aX   DTrU  G?� ^)2�h�G?���a{�X   INrV  G?���a{�X   VBrW  G?��L�x��X   JJrX  G?��L�x��X   NNSrY  G?���a{�X   VBGrZ  G?��L�x��X   JJSr[  G?��L�x��X   WRBr\  G?���a{�hMG?��L�x��X   TOr]  G?��L�x��X   CDr^  G?��L�x��X   JJRr_  G?���a{�X   VBNr`  G?���a{�X   NNra  G?��L�x��uX   NNPrb  h��rc  h h(h
c__builtin__
__main__
hNN}rd  Ntre  Rrf  �rg  Rrh  (X   INri  G?�333333X   NNSrj  G?ə�����X   RBrk  G?ə�����h�G?�333333uh�ji  �rl  h h(h
c__builtin__
__main__
hNN}rm  Ntrn  Rro  �rp  Rrq  (X   NNPrr  G?ƥjV�jWX   INrs  G?����� X   DTrt  G?�]5�]5�X   CDru  G?���X   JJrv  G?�X   NNSrw  G?�A�A�X   NNrx  G?���X   PRP$ry  G?�����h�G?��Z��Z�X   WPrz  G?�����X   VBGr{  G?����� X   ``r|  G?���� X   WDTr}  G?����� X   JJSr~  G?uPPX   PRPr  G?����� X   JJRr�  G?uPPX   VBDr�  G?uPPX   MDr�  G?uPPX   WRBr�  G?uPPX   TOr�  G?uPPuX   JJr�  ja  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   INr�  G?���4j�+X   DTr�  G?Ġ�����X   PRP$r�  G?���G���X   NNPr�  G?�;��P&X   JJr�  G?������X   VBr�  G?�=5�(>9X   WPr�  G?���&�\X   NNr�  G?���D���X   CDr�  G?{݁��vX   NNSr�  G?�݁��vh�G?�No�1�X   VBGr�  G?��݁�X   RBr�  G?���G���X   PRPr�  G?k݁��vX   VBNr�  G?`;��P%�X   WDTr�  G?k݁��vX   oovr�  G?`;��P%�NG?U��4j�+X   NNPSr�  G?k݁��vX   WRBr�  G?U��4j�+X   ``r�  G?U��4j�+uja  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   NNPr�  G?�(���X   WPr�  G?��V�AX   RBr�  G?�����X   DTr�  G?�մP#�X   PRP$r�  G?��B�YX   NNSr�  G?���|�/X   NNr�  G?�#�[EX   CDr�  G?�]~��&X   JJr�  G?���|�/X   VBGr�  G?�����X   JJSr�  G?�B�Y!dh�G?�|�.�q�X   INr�  G?���s��X   ``r�  G?��j�(�X   PRPr�  G?�*K��a�X   VBr�  G?q����X   WRBr�  G?q����uX   WPr�  j  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   PRPr�  G?�zag�zX   VBr�  G?�3s#723X   DTr�  G?ə�����X   JJr�  G?�����X   RBr�  G?�;q#�;X   CDr�  G?�����X   NNSr�  G?���ό�hMG?_����X   VBNr�  G?_����X   VBDr�  G?_����X   JJSr�  G?_����X   NNr�  G?������X   JJRr�  G?g���X   VBGr�  G?��?��X   NNPSr�  G?_����X   NNPr�  G?�����X   INr�  G?_����X   RBSr�  G?_����X   TOr�  G?_����X   PRP$r�  G?_����uj  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   VBr�  G?��q�3ʺX   RBr�  G?�2O�R��X   VBPr�  G?��ن���X   ``r�  G?w�"���uX   JJr�  j�  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   INr�  G?���S��h�G?��0=ei�X   NNr�  G?Ď��,�dX   NNSr�  G?�h�͑D�X   TOr�  G?�7]�?
X   JJr�  G?��\�t6�X   NNPr�  G?�P�XA�X   RBr�  G?��\�t6�X   VBDr�  G?q����+�X   CCr�  G?zP�XA�X   RPr�  G?q����+�X   VBNr�  G?�P�XA�X   DTr�  G?�����+�X   oovr�  G?q����+�hMG?q����+�X   WRBr�  G?q����+�uX   DTr�  j  �r�  h h(h
c__builtin__
__main__
hNN}r�  Ntr�  Rr�  �r�  Rr�  (X   JJSr�  G?�'� )*tX   NNr�  G?΍���mYX   NNPr�  G?���]��X   JJr�  G?Ռ8�_2,X   CDr�  G?��9��gX   NNSr�  G?�'� )*tX   VBNr�  G?t�9��gX   ''r�  G?t�9��gX   PRPr�  G?~��Ռ8�X   DTr�  G?���\���X   RBr�  G?��9��gX   TOr    G?��9��gh�G?~��Ռ8�X   VBr   G?t�9��guj  j�  �r   h h(h
c__builtin__
__main__
hNN}r   Ntr   Rr   �r   Rr   (X   NNr   G?�X   NNSr	   G?Ɩ�����X   JJr
   G?�X   CCr   G?�hMG?�uNh)�r   h h(h
c__builtin__
__main__
hNN}r   Ntr   Rr   �r   Rr   (X   WRBr   G?�/�A��X   INr   G?�:�c�qX   WPr   G?�c�qF:�X   NNPr   G?���!�xX   DTr   G?�A��40X   TOr   G?�F:�c�X   CDr   G?���ajzVhMG?�Z�����X   JJr   G?�s�1�8�X   NNr   G?���!�xX   VBGr   G?�c�qF:�X   VBNr   G?���	��X   RBr   G?���ajzVX   VBZr   G?r��!�xX   NNSr   G?�/�A��4X   oovr    G?{/�A��4X   VBDr!   G?���!�xX   CCr"   G?r��!�xuh)j   �r#   h h(h
c__builtin__
__main__
hNN}r$   Ntr%   Rr&   �r'   Rr(   (X   NNSr)   G?���|X   JJr*   G?�]E�t]X   VBGr+   G?�d�6M�eX   INr,   G?���|X   WPr-   G?���|X   RBr.   G?�E�t]FX   CCr/   G?���|X   NNPr0   G?�E�t]FX   PRPr1   G?�&ɲl�'X   VBZr2   G?���|NG?���|X   PRP$r3   G?�E�t]FX   VBDr4   G?���|X   DTr5   G?���|uj   j)   �r6   h h(h
c__builtin__
__main__
hNN}r7   Ntr8   Rr9   �r:   Rr;   (X   VBPr<   G?�oM�7�X   VBDr=   G?���g�Q�X   VBNr>   G?���J3�)X   CCr?   G?�B�Y!dX   TOr@   G?��`v���X   WDTrA   G?��`v���X   INrB   G?��B�YX   JJrC   G?�B�Y!dX   MDrD   G?���g�Q�X   NNrE   G?��`v���X   VBGrF   G?�B�Y!dX   RBrG   G?��`v���X   VBrH   G?��`v���X   NNPrI   G?��`v���X   DTrJ   G?��`v���X   VBZrK   G?��`v���uj<   j�  �rL   h h(h
c__builtin__
__main__
hNN}rM   NtrN   RrO   �rP   RrQ   (X   VBNrR   G?���N��X   VBDrS   G?���N��h�G?�Bd�*"yX   RPrT   G?tm�4Y`fX   INrU   G?�����mX   TOrV   G?��m�4YX   VBrW   G?ڧCL��X   VBZrX   G?���N��X   MDrY   G?�&�Q�`X   RBrZ   G?��A�o��X   VBGr[   G?�����sX   NNPr\   G?~��N��X   oovr]   G?tm�4Y`fX   NNSr^   G?tm�4Y`fX   JJr_   G?�����X   DTr`   G?�m�4Y`fX   NNra   G?�m�4Y`fX   VBPrb   G?��7���SX   NNPSrc   G?~��N��hMG?tm�4Y`fX   RBSrd   G?tm�4Y`fX   CCre   G?tm�4Y`fX   PRPrf   G?tm�4Y`fX   ``rg   G?�m�4Y`fuj�  jR   �rh   h h(h
c__builtin__
__main__
hNN}ri   Ntrj   Rrk   �rl   Rrm   (h�G?�X��Ƈ�X   INrn   G?����hX   VBNro   G?���/9X   TOrp   G?���/9X   RBSrq   G?���/9X   NNrr   G?���/9X   VBDrs   G?���/9uX   VBDrt   j�  �ru   h h(h
c__builtin__
__main__
hNN}rv   Ntrw   Rrx   �ry   Rrz   (h�G?��W��X   NNr{   G?�D=��X   INr|   G?ƫ+[��7X   NNSr}   G?�B[=t�0X   JJr~   G?�U�����X   NNPr   G?����?WX   TOr�   G?�K)ًX   WRBr�   G?p��] X   PRP$r�   G?H!-��@X   VBNr�   G?�)yh�X   CCr�   G?�W���hMG?s���TX   RBr�   G?�[�}�&X   VBGr�   G?x!-��@X   VBr�   G?p��] X   NNPSr�   G?����TX   VBZr�   G?H!-��@X   ''r�   G?b�7�X   VBDr�   G?^)yh�X   CDr�   G?p��] X   DTr�   G?e���NG?b�7�X   oovr�   G?R�7�X   JJRr�   G?X!-��@X   VBPr�   G?H!-��@X   JJSr�   G?H!-��@X   WPr�   G?R�7�X   MDr�   G?H!-��@uX   NNSr�   j�  �r�   h h(h
c__builtin__
__main__
hNN}r�   Ntr�   Rr�   �r�   Rr�   (X   VBPr�   G?f���MX   WPr�   G?t-f%��h�G?��`W�X   TOr�   G?�{���aX   INr�   G?����0~�X   NNPr�   G?{�����X   DTr�   G?v���MX   JJr�   G?�n�L�	�X   RBr�   G?�B���̤X   CCr�   G?mYNª\gX   NNSr�   G?�B���̤X   VBNr�   G?�-f%��X   RPr�   G?�mÕ&�X   PRPr�   G?]YNª\gX   VBGr�   G?����MhMG?V���MX   WDTr�   G?V���MX   WRBr�   G?f���MX   NNr�   G?����MX   ``r�   G?]YNª\gX   oovr�   G?MYNª\gX   VBDr�   G?]YNª\gX   JJSr�   G?]YNª\gX   NNPSr�   G?MYNª\gNG?MYNª\gX   VBr�   G?V���MX   VBZr�   G?V���MX   JJRr�   G?]YNª\gX   PRP$r�   G?V���MX   CDr�   G?MYNª\guj�  j�   �r�   h h(h
c__builtin__
__main__
hNN}r�   Ntr�   Rr�   �r�   Rr�   (X   NNPr�   G?�a�a�X   VBNr�   G?�a�a�X   WPr�   G?�a�a�X   NNSr�   G?�a�a�X   CCr�   G?�a�a�X   INr�   G?�I$�I$�X   TOr�   G?�a�a�ujS  j7  �r�   h h(h
c__builtin__
__main__
hNN}r�   Ntr�   Rr�   �r�   Rr�   (X   INr�   G?�      X   NNSr�   G?�      X   CCr�   G?�      X   JJr�   G?�      h�G?�      X   NNr�   G?�      X   NNPr�   G?�      X   RBr�   G?�      X   VBNr�   G?�      uX   VBGr�   j�  �r�   h h(h
c__builtin__
__main__
hNN}r�   Ntr�   Rr�   �r�   Rr�   (X   TOr�   G?�A�A�X   INr�   G?ƍh֍h�X   WPr�   G?��8�8h�G?����� X   VBNr�   G?�5�Z5�ZX   VBr�   G?��_�_X   JJr�   G?�A�A�X   RBr�   G?��K��K�X   NNPr�   G?��8�8X   NNr�   G?�a�a�X   VBZr�   G?��8�8X   CDr�   G?��8�8X   VBGr�   G?��8�8NG?��8�8X   VBDr�   G?��8�8X   DTr�   G?�a�a�X   JJRr�   G?��8�8X   VBPr�   G?��8�8X   NNSr�   G?�A�A�X   CCr�   G?��8�8uj�  j�   �r�   h h(h
c__builtin__
__main__
hNN}r�   Ntr�   Rr�   �r�   Rr�   (X   VBGr�   G?�$6Qz7SX   NNPr�   G?�%���N�X   CDr�   G?���J�iX   DTr�   G?ή�P�X   VBr�   G?�-C���(X   PRPr�   G?�$6Qz7X   PRP$r�   G?�$6Qz7Sh�G?���X	X   NNr�   G?�!1ʰX   WPr�   G?�-C���X   WRBr�   G?�-C���(X   NNSr�   G?�$6Qz7X   INr�   G?�$6Qz7X   RBr�   G?�*?_��X   WDTr�   G?�$6Qz7SX   ``r�   G?p$6Qz7X   VBNr�   G?p$6Qz7X   JJr !  G?x$6Qz7ShMG?p$6Qz7X   NNPSr!  G?p$6Qz7uj�   j�   �r!  h h(h
c__builtin__
__main__
hNN}r!  Ntr!  Rr!  �r!  Rr!  (X   PRP$r!  G?���a{�X   DTr	!  G?�B�b]X   PRPr
!  G?�-f%��X   NNPr!  G?���w͏X   NNr!  G?���w͏X   JJr!  G?�d���)�X   NNSr!  G?�{���aX   RBr!  G?�-f%��h�G?����xX   VBNr!  G?�p<�2qX   INr!  G?�-f%��X   JJRr!  G?�D8��JX   RPr!  G?�-f%��X   CCr!  G?�-f%��hMG?�D8��JX   WPr!  G?�-f%��X   VBDr!  G?�D8��JX   VBGr!  G?�-f%��X   TOr!  G?�D8��Juj�  h��r!  h h(h
c__builtin__
__main__
hNN}r!  Ntr!  Rr!  �r!  Rr!  (NG?�������X   DTr!  G?�������X   ``r !  G?�������X   NNPr!!  G?�������uX   DTr"!  j�  �r#!  h h(h
c__builtin__
__main__
hNN}r$!  Ntr%!  Rr&!  �r'!  Rr(!  (X   INr)!  G?�A�A�X   NNr*!  G?�+�+�X   ``r+!  G?��8�8X   NNSr,!  G?��y�yX   JJr-!  G?�����X   NNPr.!  G?�a�a�X   TOr/!  G?���h�G?�AAX   WPr0!  G?z��X   RBr1!  G?���X   CDr2!  G?�AAX   CCr3!  G?��8�8X   DTr4!  G?���X   ''r5!  G?z��X   oovr6!  G?z��X   WRBr7!  G?��8�8X   VBPr8!  G?z��X   NNPSr9!  G?z��uX   VBNr:!  jR  �r;!  h h(h
c__builtin__
__main__
hNN}r<!  Ntr=!  Rr>!  �r?!  Rr@!  (X   DTrA!  G?�w���X   VBrB!  G?�Z3C���X   WPrC!  G?����g��X   NNPrD!  G?���͵_�X   INrE!  G?��q���h�G?�[ғN1�X   WRBrF!  G?l�w���X   PRP$rG!  G?sw���X   JJrH!  G?��Ga��{X   PRPrI!  G?g\x�HX   NNrJ!  G?�jN�\X   WDTrK!  G?p�:�=��X   NNSrL!  G?�9�'�X   RBrM!  G?��:�=��X   TOrN!  G?_%�D#
�X   VBGrO!  G?v9�'�X   JJSrP!  G?T����#X   CDrQ!  G?_%�D#
�X   RBSrR!  G?D����#X   NNPSrS!  G?D����#NG?D����#X   VBNrT!  G?Y���r��X   oovrU!  G?O%�D#
�X   ``rV!  G?T����#X   CCrW!  G?D����#hMG?D����#uh�j�  �rX!  h h(h
c__builtin__
__main__
hNN}rY!  NtrZ!  Rr[!  �r\!  Rr]!  (X   INr^!  G?� � �X   VBNr_!  G?�A�A�X   VBZr`!  G?�A�A�X   POSra!  G?�A�A�h�G?�A�A�NG?�i�i�hMG?�A�A�X   DTrb!  G?�A�A�X   VBDrc!  G?��;�;X   TOrd!  G?�A�A�X   oovre!  G?�A�A�X   NNrf!  G?�A�A�X   MDrg!  G?�A�A�uj	  h��rh!  h h(h
c__builtin__
__main__
hNN}ri!  Ntrj!  Rrk!  �rl!  Rrm!  (X   NNSrn!  G?�`1�`X   INro!  G?�E�t]FhMG?��A)��X   NNPrp!  G?��A)��X   VBNrq!  G?���0�h�G?�E�t]FX   NNrr!  G?�E�t]FX   JJrs!  G?���0�X   CCrt!  G?��A)��X   POSru!  G?���0�X   VBGrv!  G?��A)��X   JJRrw!  G?��A)��X   CDrx!  G?���0�X   TOry!  G?��A)��X   DTrz!  G?���0�ujJ  j�  �r{!  h h(h
c__builtin__
__main__
hNN}r|!  Ntr}!  Rr~!  �r!  Rr�!  (X   NNr�!  G?�zд�TX   VBDr�!  G?�F-��DX   VBZr�!  G?�F-��DX   RBr�!  G?�[׹6�X   VBNr�!  G?ũ�g��X   PRP$r�!  G?����ǍFX   DTr�!  G?�=���aVX   NNSr�!  G?���D�RX   NNPr�!  G?�/�	uX   RBSr�!  G?xh���݅X   INr�!  G?�/�	uX   JJr�!  G?��F-�X   WPr�!  G?��+�~X   TOr�!  G?�J�s=hMG?mJ�s=X   VBGr�!  G?��+�~X   CCr�!  G?}J�s=X   JJRr�!  G?��+�~X   WRBr�!  G?�F-��DX   MDr�!  G?c�+�~X   VBPr�!  G?�F-��DX   CDr�!  G?�J�s=X   PRPr�!  G?�F-��DX   VBr�!  G?s�+�~X   oovr�!  G?�F-��DX   RPr�!  G?mJ�s=h�G?c�+�~X   ``r�!  G?�F-��Duj�  j�!  �r�!  h h(h
c__builtin__
__main__
hNN}r�!  Ntr�!  Rr�!  �r�!  Rr�!  (X   INr�!  G?�|���X   VBDr�!  G?�:'0��MX   NNPr�!  G?���읚qX   VBZr�!  G?�� ��F�h�G?���U�FX   VBNr�!  G?�,u&"��X   NNr�!  G?���<�XhMG?���읚qX   WDTr�!  G?��t�B)X   TOr�!  G?�.�k	bX   VBr�!  G?�d�ҳX   DTr�!  G?��-�ȖX   NNSr�!  G?�p�ZϿ�X   JJr�!  G?�� ��F�X   CCr�!  G?�p�ZϿ�X   RBr�!  G?��ҳ;X   VBGr�!  G?��-�ȖX   RBSr�!  G?d:'0��MX   POSr�!  G?~W:��tX   MDr�!  G?z�4@�=�X   WRBr�!  G?p� ��F�X   VBPr�!  G?d:'0��MX   PRP$r�!  G?j�4@�=�X   JJRr�!  G?Z�4@�=�X   oovr�!  G?d:'0��MNG?Z�4@�=�X   CDr�!  G?d:'0��MX   WPr�!  G?j�4@�=�X   ``r�!  G?Z�4@�=�uj  j�  �r�!  h h(h
c__builtin__
__main__
hNN}r�!  Ntr�!  Rr�!  �r�!  Rr�!  (X   DTr�!  G?�����X   PRPr�!  G?�M�l���X   TOr�!  G?����LX   WPr�!  G?�l�����X   VBGr�!  G?���]h�X   VBNr�!  G?��[���X   JJr�!  G?��M�l�X   CDr�!  G?~�|� h�G?�M�l���X   RBr�!  G?��{���X   CCr�!  G?~�|� X   NNSr�!  G?�M�l���X   NNr�!  G?�~[ i7�hMG?~�|� X   INr�!  G?�|z �w�X   oovr�!  G?v��]h�X   NNPr�!  G?���]h�X   JJRr�!  G?~�|� X   PRP$r�!  G?v��]h�X   RBSr�!  G?n�|� X   JJSr�!  G?���M�,�X   POSr�!  G?n�|� X   VBPr�!  G?n�|� X   ``r�!  G?���M�,�X   VBDr�!  G?n�|� X   RPr�!  G?n�|� uX   DTr�!  j�  �r�!  h h(h
c__builtin__
__main__
hNN}r�!  Ntr�!  Rr�!  �r�!  Rr�!  (X   VBZr�!  G?�5�yC^X   JJr�!  G?�5�yC^X   VBNr�!  G?�򆼡�(h�G?�ה5�yX   CCr�!  G?�򆼡�(X   VBPr�!  G?�򆼡�(X   VBDr�!  G?�򆼡�(uj  j�  �r�!  h h(h
c__builtin__
__main__
hNN}r�!  Ntr�!  Rr�!  �r�!  Rr�!  (X   NNr�!  G?�jt�F�X   JJr�!  G?���r5:X   PRPr�!  G?���r5:X   CDr�!  G?�jt�F�X   PRP$r�!  G?�F�eb��X   DTr�!  G?�ᕋg�X   VBNr�!  G?����[X   RBr�!  G?�ᕋg�X   NNSr�!  G?�X�~��zX   NNPr�!  G?�X�~��zX   VBGr�!  G?�jt�F�X   INr�!  G?��X�~�X   WDTr�!  G?�F�eb��X   VBPr�!  G?�F�eb��X   ``r�!  G?�F�eb��X   TOr�!  G?�jt�F�uX   WRBr�!  h@�r�!  h h(h
c__builtin__
__main__
hNN}r�!  Ntr�!  Rr "  �r"  Rr"  (X   PRPr"  G?�m�ڂX   DTr"  G?�wU�uX   NNSr"  G?�0`��X   VBr"  G?��q�-'X   NNPr"  G?�����:�X   CDr"  G?����<X   JJr	"  G?��!�X   PRP$r
"  G?sY�5�pX   oovr"  G?i�4��@X   NNr"  G?�ځ�m�X   RBr"  G?����<X   VBZr"  G?i�4��@X   JJRr"  G?i�4��@X   VBGr"  G?y�4��@X   JJSr"  G?i�4��@uX   WPr"  ji  �r"  h h(h
c__builtin__
__main__
hNN}r"  Ntr"  Rr"  �r"  Rr"  (X   NNr"  G?��m��m�X   NNSr"  G?�I$�I$�uX   NNr"  jj  �r"  h h(h
c__builtin__
__main__
hNN}r"  Ntr"  Rr"  �r "  Rr!"  (X   WDTr""  G?�X   INr#"  G?�������h�G?�X   DTr$"  G?�������X   NNr%"  G?�������X   WRBr&"  G?�X   ''r'"  G?�������X   NNPr("  G?�X   CDr)"  G?�X   PRP$r*"  G?�X   JJr+"  G?�X   RBr,"  G?�X   PRPr-"  G?�X   TOr."  G?�X   CCr/"  G?�X   VBGr0"  G?�ujj  j""  �r1"  h h(h
c__builtin__
__main__
hNN}r2"  Ntr3"  Rr4"  �r5"  Rr6"  (X   JJr7"  G?�E�t]FX   NNPr8"  G?�E�t]FX   VBDr9"  G?�E�t]FX   NNSr:"  G?�t]E�tuj�  j�  �r;"  h h(h
c__builtin__
__main__
hNN}r<"  Ntr="  Rr>"  �r?"  Rr@"  (X   INrA"  G?�
=p��
X   NNrB"  G?�333333h�G?�z�G�{X   RBrC"  G?�z�G�{X   JJrD"  G?��Q��hMG?�z�G�{X   NNSrE"  G?�z�G�{X   VBGrF"  G?�z�G�{uX   CDrG"  j-  �rH"  h h(h
c__builtin__
__main__
hNN}rI"  NtrJ"  RrK"  �rL"  RrM"  (X   NNPrN"  G?���Ol�X   CDrO"  G?���#uX   VBDrP"  G?�3�n�DX   VBGrQ"  G?v�I
�=X   DTrR"  G?���N��X   JJrS"  G?���N��X   RBrT"  G?��I
�=X   JJRrU"  G?��r+�}�X   INrV"  G?��I
�=X   oovrW"  G?����S�X   VBrX"  G?v�I
�=X   WDTrY"  G?v�I
�=X   VBPrZ"  G?v�I
�=X   WPr["  G?v�I
�=X   WRBr\"  G?v�I
�=X   NNSr]"  G?v�I
�=X   PRP$r^"  G?v�I
�=X   VBNr_"  G?����S�uj�  jO"  �r`"  h h(h
c__builtin__
__main__
hNN}ra"  Ntrb"  Rrc"  �rd"  Rre"  (hMG?�/�A��4h�G?�_�յ�}X   WPrf"  G?�*J���X   NNPrg"  G?���!�xX   NNrh"  G?��S^e1X   INri"  G?���ajzVX   RBSrj"  G?x*J���X   NNSrk"  G?�^e1�SX   JJrl"  G?�*J���X   WRBrm"  G?���!�xX   VBDrn"  G?�% �RPX   MDro"  G?x*J���X   TOrp"  G?�*J���X   VBNrq"  G?���!�xNG?�*J���X   VBPrr"  G?���!�xX   WDTrs"  G?x*J���X   RBrt"  G?���!�xX   CCru"  G?x*J���X   POSrv"  G?���!�xX   VBrw"  G?x*J���X   CDrx"  G?x*J���X   VBZry"  G?x*J���uhMjm  �rz"  h h(h
c__builtin__
__main__
hNN}r{"  Ntr|"  Rr}"  �r~"  Rr"  (X   VBZr�"  G?�������X   NNr�"  G?�������X   CDr�"  G?�������X   NNPr�"  G?�������X   VBDr�"  G?�������X   NNSr�"  G?�������X   VBPr�"  G?�������X   INr�"  G?�UUUUUUX   JJr�"  G?�X   MDr�"  G?�UUUUUUX   VBGr�"  G?�X   PRPr�"  G?�������uX   PRPr�"  j�  �r�"  h h(h
c__builtin__
__main__
hNN}r�"  Ntr�"  Rr�"  �r�"  Rr�"  (X   NNPr�"  G?�      X   VBNr�"  G?�      X   DTr�"  G?�      X   PRPr�"  G?�      X   NNSr�"  G?�      X   RBr�"  G?�      X   PRP$r�"  G?�      X   VBGr�"  G?�      X   VBDr�"  G?�      X   WPr�"  G?�      X   CCr�"  G?�      uj
  hM�r�"  h h(h
c__builtin__
__main__
hNN}r�"  Ntr�"  Rr�"  �r�"  Rr�"  (X   VBGr�"  G?��U̴�X   CCr�"  G?�����:X   NNPr�"  G?��g��k�X   WPr�"  G?����'�X   WDTr�"  G?��&��#X   WRBr�"  G?��ͣ��X   NNSr�"  G?��9Z��pX   INr�"  G?�q�q�X   JJRr�"  G?]����LX   JJr�"  G?�@��I5�X   DTr�"  G?�OEz�5X   RBr�"  G?�a�jQ"�X   NNr�"  G?�ƥ/�X   VBPr�"  G?�?jȂ��X   PRPr�"  G?z�&��#X   NNPSr�"  G?va�jQ"�X   VBNr�"  G?��qO��;X   TOr�"  G?fa�jQ"�X   ''r�"  G?m����LX   VBr�"  G?r���G�X   CDr�"  G?}����LX   JJSr�"  G?]����LX   VBDr�"  G?�?jȂ��X   VBZr�"  G?�����LX   PRP$r�"  G?fa�jQ"�X   oovr�"  G?��qO��;h�G?]����LX   ``r�"  G?]����LuhMj,  �r�"  h h(h
c__builtin__
__main__
hNN}r�"  Ntr�"  Rr�"  �r�"  Rr�"  (h�G?��_�_X   WRBr�"  G?�z�G�{X   TOr�"  G?���'EX   VBGr�"  G?�A�A�X   PRP$r�"  G?�g��4��X   CCr�"  G?�g��4��hMG?�g��4��X   DTr�"  G?�z�G�{X   WPr�"  G?�A�A�X   VBDr�"  G?�z�G�{X   INr�"  G?э�'EX   RBr�"  G?�A�A�X   VBNr�"  G?�cyj��X   VBZr�"  G?�g��4��X   NNPr�"  G?���'EX   VBPr�"  G?���'EX   WDTr�"  G?�g��4��X   NNr�"  G?�g��4��X   JJr�"  G?�g��4��X   PRPr�"  G?�g��4��X   VBr�"  G?�g��4��X   oovr�"  G?�g��4��X   CDr�"  G?�g��4��uj�	  jC  �r�"  h h(h
c__builtin__
__main__
hNN}r�"  Ntr�"  Rr�"  �r�"  Rr�"  (X   JJr�"  G?ה5�yCX   PRPr�"  G?�ה5�yX   WDTr�"  G?�򆼡�(X   VBGr�"  G?�ה5�yh�G?�5�yC^X   DTr�"  G?҆���(lX   NNSr�"  G?��5�yCX   INr�"  G?�򆼡�(X   PRP$r�"  G?�5�yC^X   NNr�"  G?�򆼡�(X   oovr�"  G?�򆼡�(X   NNPr�"  G?�5�yC^X   RBr�"  G?�5�yC^X   CDr�"  G?�򆼡�(X   VBNr�"  G?�򆼡�(X   MDr�"  G?�򆼡�(uX   VBPr�"  jH  �r�"  h h(h
c__builtin__
__main__
hNN}r�"  Ntr�"  Rr�"  �r�"  Rr�"  (X   NNSr�"  G?�0_}T~�X   NNr�"  G?�y��hH�X   INr�"  G?�mOxM�>h�G?��MEkX   TOr�"  G?� �I��)X   CCr�"  G?�)&�y?X   JJr�"  G?���=��X   NNPr�"  G?����"<�X   VBGr�"  G?��MEkhMG?�ؼw\��X   VBNr�"  G?�'��-�1X   NNPSr�"  G?tb�s�!X   VBr #  G?� �I��)X   WPr#  G?db�s�!X   VBZr#  G?^'��-�1X   PRPr#  G?^'��-�1X   RBr#  G?�����e%X   WRBr#  G?i �I��)X   ''r#  G?^'��-�1X   ``r#  G?Tb�s�!X   DTr#  G?v����e%X   CDr	#  G?db�s�!X   VBDr
#  G?db�s�!X   VBPr#  G?Tb�s�!X   oovr#  G?db�s�!NG?Tb�s�!X   RBSr#  G?^'��-�1X   JJRr#  G?Tb�s�!X   POSr#  G?^'��-�1uX   WRBr#  hA�r#  h h(h
c__builtin__
__main__
hNN}r#  Ntr#  Rr#  �r#  Rr#  (X   NNPr#  G?�kጹO�X   PRPr#  G?���϶�VX   VBNr#  G?���eX   DTr#  G?�Wo�sGX   VBr#  G?����y�mX   NNr#  G?�E�t]FX   JJr#  G?�J�m/�
X   oovr#  G?{��F�X   JJSr#  G?{��F�X   RBr #  G?������X   VBGr!#  G?�Q�����X   VBZr"#  G?[��F�X   RBSr##  G?d�U�.X   INr$#  G?k��F�X   CDr%#  G?����@�X   VBDr&#  G?K��F�X   ``r'#  G?t�U�.X   NNSr(#  G?h\8���X   PRP$r)#  G?k��F�X   TOr*#  G?K��F�uX   RBr+#  j�  �r,#  h h(h
c__builtin__
__main__
hNN}r-#  Ntr.#  Rr/#  �r0#  Rr1#  (h�G?Ԫ�����X   VBDr2#  G?�UUUUUUX   WRBr3#  G?�UUUUUUX   NNr4#  G?�      X   VBPr5#  G?�UUUUUUX   TOr6#  G?�      X   VBZr7#  G?�UUUUUUX   JJr8#  G?�      X   INr9#  G?�      X   VBr:#  G?�UUUUUUX   MDr;#  G?�UUUUUUuX   VBPr<#  j
  �r=#  h h(h
c__builtin__
__main__
hNN}r>#  Ntr?#  Rr@#  �rA#  RrB#  (X   NNPrC#  G?�v��!gX   INrD#  G?�q�q�X   VBNrE#  G?�6���nX   TOrF#  G?����� X   NNrG#  G?��fA�h�G?��fA�X   JJrH#  G?��
�
X   PRP$rI#  G?l��X   WPrJ#  G?�a&a&X   RBrK#  G?�A�A�X   CDrL#  G?r��h*�X   NNSrM#  G?�,k�b�X   DTrN#  G?��fA�hMG?�VZ�fX   JJRrO#  G?b��h*�X   RPrP#  G?�VZ�fX   JJSrQ#  G?b��h*�X   CCrR#  G?~W:��tX   WRBrS#  G?�֒��=iX   RBSrT#  G?b��h*�X   VBGrU#  G?l��X   WDTrV#  G?R��h*�X   VBDrW#  G?R��h*�X   PRPrX#  G?gV��umNG?R��h*�X   VBrY#  G?R��h*�X   oovrZ#  G?l��X   ``r[#  G?gV��umX   ''r\#  G?R��h*�X   VBPr]#  G?R��h*�ujx  j  �r^#  h h(h
c__builtin__
__main__
hNN}r_#  Ntr`#  Rra#  �rb#  Rrc#  (X   VBNrd#  G?��j���X   VBre#  G?�BG�X�X   DTrf#  G?�$��6X   WRBrg#  G?|�Y$�ѻX   RBrh#  G?�^%� �X   oovri#  G?�K��eyX   VBGrj#  G?�$��6X   NNPrk#  G?�$��6X   INrl#  G?��Y$�ѻX   CDrm#  G?�&h�ɱ
h�G?����SnX   WPrn#  G?�K��eyX   JJro#  G?�}h݅r�X   NNrp#  G?�$��6X   VBPrq#  G?q&h�ɱ
X   TOrr#  G?��W��X   JJRrs#  G?�&h�ɱ
X   ``rt#  G?f���bAbX   CCru#  G?a&h�ɱ
X   PRP$rv#  G?a&h�ɱ
X   PRPrw#  G?a&h�ɱ
hMG?l�Y$�ѻX   NNPSrx#  G?V���bAbX   RPry#  G?a&h�ɱ
X   VBZrz#  G?a&h�ɱ
X   NNSr{#  G?a&h�ɱ
X   VBDr|#  G?a&h�ɱ
uX   VBZr}#  j�!  �r~#  h h(h
c__builtin__
__main__
hNN}r#  Ntr�#  Rr�#  �r�#  Rr�#  (X   NNPr�#  G?�      X   RBr�#  G?�ډ]���X   JJRr�#  G?������X   JJr�#  G?�ډ]���X   DTr�#  G?Ԯ�J�D�X   INr�#  G?��Q+��X   NNr�#  G?��Q+��X   WPr�#  G?������X   VBGr�#  G?��Q+��X   VBNr�#  G?�81�8X   VBr�#  G?��Q+��X   PRPr�#  G?������X   CDr�#  G?������X   CCr�#  G?������X   WRBr�#  G?������ujc  j  �r�#  h h(h
c__builtin__
__main__
hNN}r�#  Ntr�#  Rr�#  �r�#  Rr�#  (X   NNSr�#  G?��Gq�wX   NNr�#  G?��'���{X   INr�#  G?��Cy�8X   TOr�#  G?��WQ]Eh�G?�Cy�7�X   NNPr�#  G?��o!��X   JJr�#  G?��/���X   VBNr�#  G?��Gq�wX   VBGr�#  G?��[Im%�X   WPr�#  G?c�Oa=��X   RBr�#  G?��k)���X   VBr�#  G?�Ki-���X   CCr�#  G?�[Im%��X   POSr�#  G?c�Oa=��X   DTr�#  G?��w�GqhMG?��g1��sX   ''r�#  G?k�o!���X   RBSr�#  G?c�Oa=��X   WRBr�#  G?g�_A}�X   CDr�#  G?o���X   oovr�#  G?o���X   RPr�#  G?O���X   NNPSr�#  G?k�o!���X   VBDr�#  G?O���X   VBZr�#  G?g�_A}�X   JJRr�#  G?_���NG?c�Oa=��X   WDTr�#  G?W�_A}�X   PRPr�#  G?W�_A}�X   JJSr�#  G?O���X   ``r�#  G?O���uhMj�"  �r�#  h h(h
c__builtin__
__main__
hNN}r�#  Ntr�#  Rr�#  �r�#  Rr�#  (X   WPr�#  G?�h�i?�X   JJr�#  G?���.K-�X   NNSr�#  G?�]�;Y�PX   NNPr�#  G?�D���1X   MDr�#  G?�����X   DTr�#  G?��{s$�X   NNr�#  G?� ʕ�k�X   INr�#  G?�}O"ljX   VBZr�#  G?�����X   VBr�#  G?��^���=X   VBDr�#  G?�ț��fX   RBr�#  G?��^���=X   VBGr�#  G?�}O"ljX   CDr�#  G?�}O"ljX   ``r�#  G?r����X   JJSr�#  G?�^���=X   PRPr�#  G?yR�s�X   VBNr�#  G?yR�s�X   VBPr�#  G?�����X   JJRr�#  G?yR�s�X   TOr�#  G?yR�s�X   oovr�#  G?r����X   WDTr�#  G?iR�s�X   WRBr�#  G?�^���=X   PRP$r�#  G?iR�s�X   NNPSr�#  G?r����uj�"  j�#  �r�#  h h(h
c__builtin__
__main__
hNN}r�#  Ntr�#  Rr�#  �r�#  Rr�#  (X   JJr�#  G?����h�G?ʡ���a�X   INr�#  G?�}l=�3�X   NNr�#  G?����X   RBr�#  G?��[wX   VBZr�#  G?��.c��X   WDTr�#  G?{}l=�3�X   VBDr�#  G?�.c��`7X   NNPr�#  G?�}l=�3�X   MDr�#  G?��.c��X   VBPr�#  G?�.c��`7X   NNSr�#  G?{}l=�3�X   CDr�#  G?{}l=�3�X   TOr�#  G?��.c��X   VBr�#  G?{}l=�3�uX   VBr�#  j�  �r�#  h h(h
c__builtin__
__main__
hNN}r�#  Ntr�#  Rr�#  �r�#  Rr�#  (h�G?�E�t]X   INr�#  G?�t]E�tX   TOr�#  G?�E�t]X   VBr�#  G?����`jX   VBPr�#  G?�]E�t]X   WDTr�#  G?�t]E�tX   CCr�#  G?��m��m�hMG?���B~VqX   DTr�#  G?s�O��X   VBZr�#  G?j��`jc�X   VBNr�#  G?��Lw�X   POSr�#  G?wE�t]FX   PRPr�#  G?c�O��X   RBr�#  G?�B~Vq	�X   WPr�#  G?z��`jc�X   VBGr�#  G?��B~Vq
X   NNr�#  G?����B~VX   JJr�#  G?�E�t]FNG?j��`jc�X   RPr $  G?Z��`jc�X   VBDr$  G?j��`jc�X   JJRr$  G?j��`jc�X   CDr$  G?c�O��X   NNPr$  G?Z��`jc�X   WRBr$  G?s�O��X   MDr$  G?j��`jc�X   NNSr$  G?}�Lw�5X   oovr$  G?Z��`jc�uj}  j�  �r	$  h h(h
c__builtin__
__main__
hNN}r
$  Ntr$  Rr$  �r$  Rr$  (X   VBNr$  G?��az�DTX   INr$  G?�ƚ�'-X   VBDr$  G?�f	=�X   POSr$  G?�8{�}��X   CCr$  G?�',��[X   RBr$  G?�',��[h�G?�ڥ���X   NNr$  G?���n< �X   NNPr$  G?�OB�]�X   DTr$  G?}',��[X   ''r$  G?�',��[X   VBPr$  G?��az�DTX   NNSr$  G?��az�DThMG?��G|ϷX   VBZr$  G?��G|ϷX   VBGr$  G?��az�DTX   TOr$  G?�',��[X   CDr$  G?��az�DTX   WRBr$  G?}',��[X   NNPSr $  G?��az�DTX   MDr!$  G?}',��[X   VBr"$  G?�',��[X   JJr#$  G?�8{�}��X   oovr$$  G?}',��[uj$  j�  �r%$  h h(h
c__builtin__
__main__
hNN}r&$  Ntr'$  Rr($  �r)$  Rr*$  (X   INr+$  G?�q�q�X   VBNr,$  G?�X   JJr-$  G?��l�lX   NNr.$  G?�X   TOr/$  G?�X   PRPr0$  G?�X   NNSr1$  G?��l�lX   DTr2$  G?�X   WRBr3$  G?��l�lX   RPr4$  G?��l�lh�G?�X   JJRr5$  G?��l�lX   WPr6$  G?��l�luj�  jD  �r7$  h h(h
c__builtin__
__main__
hNN}r8$  Ntr9$  Rr:$  �r;$  Rr<$  (X   RBr=$  G?�%���N�X   VBDr>$  G?˩~=\
X   VBr?$  G?�$6Qz7X   NNr@$  G?�$6Qz7X   MDrA$  G?p$6Qz7X   DTrB$  G?��y���X   VBNrC$  G?��y���X   INrD$  G?�%���N�X   TOrE$  G?�!1ʰh�G?�-C���X   VBPrF$  G?�$6Qz7X   ``rG$  G?p$6Qz7X   WRBrH$  G?�$6Qz7X   VBZrI$  G?�-C���X   VBGrJ$  G?�$6Qz7X   JJRrK$  G?�-C���X   JJrL$  G?��y���X   oovrM$  G?�*?_��X   CCrN$  G?x$6Qz7SX   NNPrO$  G?�$6Qz7X   JJSrP$  G?p$6Qz7hMG?x$6Qz7SX   RPrQ$  G?x$6Qz7SX   WDTrR$  G?p$6Qz7ujD  j=$  �rS$  h h(h
c__builtin__
__main__
hNN}rT$  NtrU$  RrV$  �rW$  RrX$  (X   VBGrY$  G?� �I��)X   INrZ$  G?�F�¿�|X   VBr[$  G?�������h�G?�i:E�X   MDr\$  G?�ؼw\��X   VBDr]$  G?��$i:X   VBPr^$  G?�j�+���X   VBNr_$  G?� �I��)X   VBZr`$  G?� �I��)X   NNra$  G?�ؼw\��X   oovrb$  G?� �I��)X   JJrc$  G?�ؼw\��X   CCrd$  G?� �I��)hMG?� �I��)X   WPre$  G?� �I��)X   TOrf$  G?�i:E�X   RBrg$  G?�i:E�X   DTrh$  G?� �I��)X   CDri$  G?�ؼw\��X   ``rj$  G?� �I��)uj=$  jY$  �rk$  h h(h
c__builtin__
__main__
hNN}rl$  Ntrm$  Rrn$  �ro$  Rrp$  (h�G?�T�+���X   RBrq$  G?�#�J+�X   INrr$  G?ļ6;��X   NNrs$  G?�#�J+�hMG?�#�J+�X   VBNrt$  G?�#�J+�X   JJru$  G?��f�宧X   NNSrv$  G?��6;��X   TOrw$  G?�T�+���X   PRP$rx$  G?���YR$�X   DTry$  G?��f�宧X   PRPrz$  G?�T�+���X   VBGr{$  G?�#�J+�X   NNPr|$  G?��6;��X   RPr}$  G?�#�J+�X   CCr~$  G?y�/���X   WPr$  G?�T�+���X   oovr�$  G?�#�J+�X   CDr�$  G?y�/���X   VBr�$  G?y�/���X   VBDr�$  G?y�/���uje#  j  �r�$  h h(h
c__builtin__
__main__
hNN}r�$  Ntr�$  Rr�$  �r�$  Rr�$  (X   NNr�$  G?���Q�X   JJr�$  G?���Q�X   CDr�$  G?��Q��X   VBDr�$  G?�z�G�{X   NNSr�$  G?��Q��X   VBZr�$  G?�z�G�{X   VBPr�$  G?��Q��uX   VBZr�$  jF  �r�$  h h(h
c__builtin__
__main__
hNN}r�$  Ntr�$  Rr�$  �r�$  Rr�$  (h�G?َ�����X   VBDr�$  G?{}l=�3�X   CDr�$  G?�.c��`7X   NNr�$  G?�1�T0}X   JJr�$  G?��ŕy�X   INr�$  G?�ŕy��RhMG?{}l=�3�X   WPr�$  G?{}l=�3�X   NNPr�$  G?{}l=�3�X   VBGr�$  G?�.c��`7X   NNSr�$  G?����X   VBZr�$  G?����X   TOr�$  G?��.c��X   VBr�$  G?��.c��uX   NNPr�$  j	  �r�$  h h(h
c__builtin__
__main__
hNN}r�$  Ntr�$  Rr�$  �r�$  Rr�$  (X   VBDr�$  G?�鮚鮛X   NNPr�$  G?����� X   VBZr�$  G?�9Ü9ÜX   CDr�$  G?�a&a&X   NNr�$  G?����� X   MDr�$  G?�a&a&X   RBr�$  G?�A�A�X   NNSr�$  G?����� X   DTr�$  G?����� X   VBPr�$  G?����� uX   TOr�$  j  �r�$  h h(h
c__builtin__
__main__
hNN}r�$  Ntr�$  Rr�$  �r�$  Rr�$  (X   NNSr�$  G?� 6@l��X   NNr�$  G?�3��P��X   NNPr�$  G?�X(�Q`�h�G?�X(�Q`�X   INr�$  G?�b�pu��X   VBr�$  G?����Zk`X   JJr�$  G?�y�HU�X   CCr�$  G?����Zk`X   NNPSr�$  G?ry�HU�X   TOr�$  G?{ 6@l��X   DTr�$  G?ry�HU�X   VBGr�$  G?ry�HU�hMG?ry�HU�X   oovr�$  G?ry�HU�uX   JJSr�$  j�  �r�$  h h(h
c__builtin__
__main__
hNN}r�$  Ntr�$  Rr�$  �r�$  Rr�$  (X   PRP$r�$  G?��C���X   DTr�$  G?��k[X   NNPr�$  G?ȸ6.��X   NNr�$  G?����pX   WPr�$  G?��kZ�X   PRPr�$  G?�����/hX   INr�$  G?��kZ�X   VBGr�$  G?�AAh�G?�AAX   WDTr�$  G?��kZ�X   JJr�$  G?����pX   VBNr�$  G?u�kZ�X   NNSr�$  G?�AAX   VBZr�$  G?u�kZ�X   CDr�$  G?�AAX   oovr�$  G?u�kZ�uj�"  jH  �r�$  h h(h
c__builtin__
__main__
hNN}r�$  Ntr�$  Rr�$  �r�$  Rr�$  (X   NNSr�$  G?�      X   NNr�$  G?�������X   JJr�$  G?�q�q�X   VBDr�$  G?uUUUUUUX   VBZr�$  G?uUUUUUUX   VBGr�$  G?lq�q�X   VBPr�$  G?|q�q�X   NNPr�$  G?�q�q�X   NNPSr�$  G?lq�q�X   RBr�$  G?lq�q�X   INr�$  G?lq�q�uX   VBPr�$  j0  �r�$  h h(h
c__builtin__
__main__
hNN}r�$  Ntr�$  Rr�$  �r�$  Rr�$  (X   INr�$  G?�9	H��h�G?��x�d��X   NNPr�$  G?�.l�O��X   DTr�$  G?�:\و�,X   VBGr�$  G?��K�1�X   WPr�$  G?�9	H��X   JJr�$  G?��K�1�X   NNr�$  G?��K�1�X   PRP$r�$  G?�Ս�n�X   JJRr�$  G?�Ս�n�X   JJSr�$  G?�9	H��X   WRBr %  G?�Ս�n�X   WDTr%  G?�9	H��NG?�9	H��X   oovr%  G?�9	H��X   TOr%  G?�Ս�n�X   RBr%  G?�Ս�n�X   VBNr%  G?�9	H��X   NNSr%  G?�Ս�n�X   CDr%  G?�9	H��uX   CDr%  j�
  �r	%  h h(h
c__builtin__
__main__
hNN}r
%  Ntr%  Rr%  �r%  Rr%  (X   VBNr%  G?�������X   NNPr%  G?�]����)X   NNr%  G?���a{�X   ``r%  G?|?����X   INr%  G?�k�Q6�%h�G?�ż�[�X   DTr%  G?ȷ�!�y�X   WDTr%  G?�/�AR��X   JJRr%  G?�/�AR��X   WPr%  G?�/�AR��X   WRBr%  G?���!�y�X   NNSr%  G?�{���aX   TOr%  G?�ż�[�X   PRP$r%  G?���a{�X   VBGr%  G?�/�AR��X   RPr%  G?�/�AR��X   VBr%  G?�/�AR��X   CDr%  G?�?����X   JJr %  G?�?����X   RBSr!%  G?|?����X   RBr"%  G?�?����X   PRPr#%  G?���a{�X   CCr$%  G?|?����X   VBDr%%  G?|?����hMG?|?����ujk  j�  �r&%  h h(h
c__builtin__
__main__
hNN}r'%  Ntr(%  Rr)%  �r*%  Rr+%  (X   ``r,%  G?�������X   NNr-%  G?�      X   JJr.%  G?�������X   NNSr/%  G?�333333X   NNPr0%  G?�������X   JJSr1%  G?�      X   CCr2%  G?�������X   VBGr3%  G?�333333h�G?�������X   RBSr4%  G?�333333X   INr5%  G?�������X   VBDr6%  G?�333333uj�  j,%  �r7%  h h(h
c__builtin__
__main__
hNN}r8%  Ntr9%  Rr:%  �r;%  Rr<%  (X   JJr=%  G?�{���aX   NNPr>%  G?�{���aX   JJSr?%  G?���a{�X   DTr@%  G?���a{�X   VBZrA%  G?���a{�X   VBNrB%  G?���a|X   VBGrC%  G?���a{�h�G?���a{�X   NNrD%  G?���a{�X   INrE%  G?�{���aujZ  j.  �rF%  h h(h
c__builtin__
__main__
hNN}rG%  NtrH%  RrI%  �rJ%  RrK%  (X   ''rL%  G?�I$�I$�h�G?�      X   VBPrM%  G?�I$�I$�X   VBDrN%  G?�m��m��X   TOrO%  G?�I$�I$�X   NNrP%  G?�I$�I$�X   INrQ%  G?�I$�I$�X   NNPSrR%  G?�m��m��uj$  hĆrS%  h h(h
c__builtin__
__main__
hNN}rT%  NtrU%  RrV%  �rW%  RrX%  (h�G?ٙ�����X   INrY%  G?��z�zX   oovrZ%  G?�PPX   NNr[%  G?�鮚鮛X   ``r\%  G?�PPX   VBGr]%  G?�PPX   TOr^%  G?�PPX   VBZr_%  G?��z�zX   JJr`%  G?�PPX   NNSra%  G?����� X   VBDrb%  G?����� hMG?����� X   MDrc%  G?�PPX   NNPrd%  G?�PPX   RBre%  G?�PPuX   PRP$rf%  h��rg%  h h(h
c__builtin__
__main__
hNN}rh%  Ntri%  Rrj%  �rk%  Rrl%  NG?�      sX   POSrm%  jT  �rn%  h h(h
c__builtin__
__main__
hNN}ro%  Ntrp%  Rrq%  �rr%  Rrs%  (X   JJrt%  G?�^rT�>#X   NNru%  G?㒤	�^X   NNSrv%  G?�{q�j�h�G?��CV��X   VBNrw%  G?��,��X   RBrx%  G?�����X   CCry%  G?�����X   VBGrz%  G?��CV��X   NNPr{%  G?���Q0�YX   ``r|%  G?z��Q0�YX   WPr}%  G?z��Q0�YuX   TOr~%  j  �r%  h h(h
c__builtin__
__main__
hNN}r�%  Ntr�%  Rr�%  �r�%  Rr�%  (X   VBr�%  G?�      X   NNPr�%  G?�      X   JJr�%  G?�      X   DTr�%  G?�      X   NNSr�%  G?�      X   PRP$r�%  G?�      uj7  jQ  �r�%  h h(h
c__builtin__
__main__
hNN}r�%  Ntr�%  Rr�%  �r�%  Rr�%  (X   CCr�%  G?|鶃P�h�G?�칆S�X   NNr�%  G?�X   INr�%  G?�}�J�~X   DTr�%  G?�I|��IX   VBGr�%  G?�I|��IX   JJr�%  G?�_+�Œ_X   NNPr�%  G?�鶃P�X   CDr�%  G?��H�|�X   VBPr�%  G?�Fy��FX   TOr�%  G?�鶃P�X   WRBr�%  G?|鶃P�X   oovr�%  G?�X   WPr�%  G?�X   VBNr�%  G?��K��X   RBr�%  G?�Fy��FX   NNSr�%  G?�Fy��FX   RPr�%  G?sFy��FhMG?|鶃P�X   VBZr�%  G?�鶃P�X   JJRr�%  G?sFy��FX   PRP$r�%  G?sFy��FX   VBDr�%  G?�ݪwD�NG?sFy��FX   VBr�%  G?�ݪwD�ujQ  j�%  �r�%  h h(h
c__builtin__
__main__
hNN}r�%  Ntr�%  Rr�%  �r�%  Rr�%  (X   VBr�%  G?�ה5�yX   RBr�%  G?�5�yC^X   JJr�%  G?�򆼡�(X   MDr�%  G?�5�yC^X   JJRr�%  G?�򆼡�(X   NNSr�%  G?�򆼡�(X   VBZr�%  G?�򆼡�(X   NNr�%  G?�򆼡�(X   INr�%  G?�5�yC^X   VBNr�%  G?�5�yC^X   VBGr�%  G?�5�yC^X   oovr�%  G?�򆼡�(X   NNPr�%  G?�򆼡�(X   VBDr�%  G?�򆼡�(X   WPr�%  G?�򆼡�(uj�  j�  �r�%  h h(h
c__builtin__
__main__
hNN}r�%  Ntr�%  Rr�%  �r�%  Rr�%  (X   VBDr�%  G?�UUUUUUX   VBPr�%  G?�      X   DTr�%  G?�UUUUUUX   VBZr�%  G?�UUUUUUX   NNr�%  G?�q�q�X   JJr�%  G?�q�q�X   MDr�%  G?�UUUUUUX   NNSr�%  G?�q�q�uj�%  j�  �r�%  h h(h
c__builtin__
__main__
hNN}r�%  Ntr�%  Rr�%  �r�%  Rr�%  (h�G?�      X   NNPr�%  G?�      NG?�������X   INr�%  G?�������X   DTr�%  G?ə�����X   NNSr�%  G?�������uX   VBNr�%  jg  �r�%  h h(h
c__builtin__
__main__
hNN}r�%  Ntr�%  Rr�%  �r�%  Rr�%  (X   JJr�%  G?���|X   NNPr�%  G?���|X   VBDr�%  G?�&ɲl�'X   VBZr�%  G?�d�6M�eX   MDr�%  G?�E�t]FX   NNr�%  G?�d�6M�eX   VBPr�%  G?���|uX   VBGr�%  j:  �r�%  h h(h
c__builtin__
__main__
hNN}r�%  Ntr�%  Rr�%  �r�%  Rr�%  (X   PRPr�%  G?�������X   VBDr�%  G?�������X   NNr�%  G?�������X   NNPr�%  G?�      X   DTr�%  G?�333333X   INr�%  G?�333333X   JJr�%  G?�������X   VBNr�%  G?�������X   VBr�%  G?�������h�G?�      X   TOr�%  G?�������uj�!  jA$  �r�%  h h(h
c__builtin__
__main__
hNN}r�%  Ntr�%  Rr�%  �r�%  Rr�%  (X   VBr�%  G?�z�G�X   INr�%  G?�z�G�{X   RBr�%  G?˅�Q�X   VBNr�%  G?��Q��X   TOr�%  G?��Q��X   VBDr�%  G?�z�G�{X   NNr�%  G?��Q��h�G?�z�G�{X   CDr &  G?�z�G�{uj	  j�  �r&  h h(h
c__builtin__
__main__
hNN}r&  Ntr&  Rr&  �r&  Rr&  (h�G?�333333X   NNr&  G?ə�����X   TOr&  G?ə�����X   CCr	&  G?�333333uj;  j�  �r
&  h h(h
c__builtin__
__main__
hNN}r&  Ntr&  Rr&  �r&  Rr&  X   VBr&  G?�      sj�	  j�  �r&  h h(h
c__builtin__
__main__
hNN}r&  Ntr&  Rr&  �r&  Rr&  (X   JJr&  G?�aq�X   NNr&  G?�_�%��`X   NNPr&  G?�B�!BX   INr&  G?��!B�X   WPr&  G?�aq�X   NNSr&  G?���,��X   ``r&  G?���=�X   VBZr&  G?jm��mX   NNPSr&  G?�x�W�yX   VBNr &  G?jm��mX   CDr!&  G?�x�W�yX   VBr"&  G?jm��mX   JJRr#&  G?jm��mX   VBGr$&  G?s��=�X   oovr%&  G?jm��mX   VBDr&&  G?jm��mh�G?s��=�X   VBPr'&  G?s��=�X   RBr(&  G?s��=�X   JJSr)&  G?s��=�ujB$  h��r*&  h h(h
c__builtin__
__main__
hNN}r+&  Ntr,&  Rr-&  �r.&  Rr/&  (X   ''r0&  G?��L�x��NG?�lߡ���X   CDr1&  G?���a{�X   ``r2&  G?��L�x��ujR  j�  �r3&  h h(h
c__builtin__
__main__
hNN}r4&  Ntr5&  Rr6&  �r7&  Rr8&  (X   JJr9&  G?�'��-�sX   WPr:&  G?����M߀X   oovr;&  G?x���JX   VBGr<&  G?�+:�ޕ X   VBNr=&  G?�4���=�X   VBr>&  G?�n��4m%X   NNr?&  G?��A�}eX   VBDr@&  G?�+:�ޕ X   RBrA&  G?�e,t��7X   NNPrB&  G?�v	2�:@X   DTrC&  G?���l֜\X   NNSrD&  G?�n��4m%X   VBPrE&  G?}n��4m%X   INrF&  G?��Z"�nX   VBZrG&  G?x���JX   NNPSrH&  G?mn��4m%X   JJRrI&  G?s�Z"�nX   JJSrJ&  G?mn��4m%X   RBSrK&  G?c�Z"�nX   MDrL&  G?mn��4m%X   WDTrM&  G?c�Z"�nX   PRP$rN&  G?c�Z"�nuj�  j9&  �rO&  h h(h
c__builtin__
__main__
hNN}rP&  NtrQ&  RrR&  �rS&  RrT&  (h�G?�:�p�~X   NNrU&  G?�}9ۊ�X   NNSrV&  G?���L1X   RBrW&  G?|�Rm_�X   INrX&  G?��3�[�&X   NNPrY&  G?� ���_X   DTrZ&  G?v1#�g�hMG?�򆼡�(X   WPr[&  G?i\��w�X   VBNr\&  G?����U�X   JJr]&  G?�S8E�aX   CCr^&  G?�1#�g�X   TOr_&  G?���[%@3X   CDr`&  G?|�Rm_�X   VBPra&  G?v1#�g�X   VBDrb&  G?o����U�X   VBrc&  G?Y\��w�X   NNPSrd&  G?Y\��w�X   VBGre&  G?i\��w�X   oovrf&  G?Y\��w�X   VBZrg&  G?Y\��w�uX   NNrh&  j  �ri&  h h(h
c__builtin__
__main__
hNN}rj&  Ntrk&  Rrl&  �rm&  Rrn&  (X   NNro&  G?�Z�����X   NNSrp&  G?�c�qF:�X   VBZrq&  G?�c�qF:�X   JJrr&  G?�Ұ�=+X   INrs&  G?�A��40X   oovrt&  G?���!�xNG?���!�xX   ``ru&  G?�/�A��4X   VBDrv&  G?�/�A��4X   CCrw&  G?��Q���X   VBPrx&  G?���!�xh�G?���ajzVX   NNPry&  G?�/�A��4X   RBrz&  G?�c�qF:�hMG?�/�A��4X   VBGr{&  G?���ajzVX   WPr|&  G?���ajzVX   MDr}&  G?���!�xX   CDr~&  G?���!�xX   DTr&  G?���ajzVX   WDTr�&  G?���!�xX   PRPr�&  G?�/�A��4X   PRP$r�&  G?���!�xuX   VBPr�&  j
  �r�&  h h(h
c__builtin__
__main__
hNN}r�&  Ntr�&  Rr�&  �r�&  Rr�&  (X   PRP$r�&  G?�[_u'X   WPr�&  G?�[_u'X   RBr�&  G?���/��X   VBNr�&  G?�[_u'h�G?���/��X   INr�&  G?����Rp�X   JJr�&  G?���/��X   NNSr�&  G?��I�A�X   NNr�&  G?�4[_uX   NNPr�&  G?���/��X   VBr�&  G?����8h#X   DTr�&  G?���/��hMG?���/��X   ''r�&  G?�[_u'X   PRPr�&  G?�[_u'X   WRBr�&  G?�[_u'X   oovr�&  G?�[_u'X   RPr�&  G?�[_u'X   VBGr�&  G?�[_u'uX   RBr�&  jf#  �r�&  h h(h
c__builtin__
__main__
hNN}r�&  Ntr�&  Rr�&  �r�&  Rr�&  (X   NNr�&  G?۴%�	{BX   JJr�&  G?�8�8�X   NNPr�&  G?�����/hX   VBNr�&  G?r����/hX   RBSr�&  G?�����/X   JJSr�&  G?���%�	{X   NNPSr�&  G?�����/hX   NNSr�&  G?�B^З�&X   VBGr�&  G?r����/hX   MDr�&  G?r����/hh�G?r����/hX   oovr�&  G?r����/hX   INr�&  G?�З�%�	X   JJRr�&  G?|q�q�X   VBDr�&  G?r����/hX   WPr�&  G?|q�q�X   RBr�&  G?|q�q�X   CDr�&  G?r����/hX   ``r�&  G?r����/huX   VBZr�&  j�  �r�&  h h(h
c__builtin__
__main__
hNN}r�&  Ntr�&  Rr�&  �r�&  Rr�&  (h�G?�X   NNr�&  G?�""""""X   JJr�&  G?љ�����X   INr�&  G?�X   NNSr�&  G?�DDDDDDX   RBr�&  G?�������X   NNPr�&  G?�X   VBNr�&  G?�������X   ''r�&  G?�������X   JJSr�&  G?�uj>  j�  �r�&  h h(h
c__builtin__
__main__
hNN}r�&  Ntr�&  Rr�&  �r�&  Rr�&  (X   JJSr�&  G?�UUUUUUX   INr�&  G?�UUUUUUX   NNSr�&  G?�UUUUUUuX   WRBr�&  jH  �r�&  h h(h
c__builtin__
__main__
hNN}r�&  Ntr�&  Rr�&  �r�&  Rr�&  (X   TOr�&  G?�rb
��X   VBGr�&  G?�Ɉ+�WX   NNPr�&  G?�l���RX   NNSr�&  G?�W& �LAh�G?�W& �LAX   DTr�&  G?�F�����X   INr�&  G?��;�6xX   JJRr�&  G?�W& �LAX   WDTr�&  G?�Ɉ+�WX   PRP$r�&  G?���1rbX   NNr�&  G?����1rX   WPr�&  G?�Ɉ+�WX   ``r�&  G?�Ɉ+�WX   PRPr�&  G?�Ɉ+�WX   JJr�&  G?�;�6w�mX   WRBr�&  G?�Ɉ+�WX   RBr�&  G?�Ɉ+�WX   VBNr�&  G?�Ɉ+�WX   VBDr�&  G?�Ɉ+�WX   oovr�&  G?�Ɉ+�WujH  j�&  �r�&  h h(h
c__builtin__
__main__
hNN}r�&  Ntr�&  Rr�&  �r�&  Rr�&  (X   NNPr�&  G?�F`F`X   WDTr�&  G?q��X   PRPr�&  G?u�^�^X   WPr�&  G?�Y��Y��X   NNr�&  G?��L��L�X   VBr�&  G?�v'bv'bX   PRP$r�&  G?���h�G?�A�A�X   DTr�&  G?�����	X   CDr�&  G?u�^�^X   JJr�&  G?�������X   NNSr�&  G?���X   NNPSr�&  G?zA�A�X   INr�&  G?���X   JJSr�&  G?jA�A�X   oovr�&  G?a��X   VBGr�&  G?jA�A�X   WRBr�&  G?jA�A�X   RBr�&  G?q��X   JJRr�&  G?jA�A�uX   DTr '  j�  �r'  h h(h
c__builtin__
__main__
hNN}r'  Ntr'  Rr'  �r'  Rr'  (X   VBNr'  G?�sL6���X   JJr'  G?���u@}X   oovr	'  G?�����i�X   CDr
'  G?�U�sX   NNPr'  G?�����i�X   NNr'  G?�sL6���X   CCr'  G?�sL6���X   INr'  G?�De�JBqX   NNSr'  G?�sL6���X   RBr'  G?�De�JBqh�G?�De�JBquj�  j'  �r'  h h(h
c__builtin__
__main__
hNN}r'  Ntr'  Rr'  �r'  Rr'  (h�G?ӱ;�;X   INr'  G?�UUUUUUX   DTr'  G?�A�A�X   TOr'  G?�A�A�X   NNSr'  G?�A�A�X   JJr'  G?�A�A�uX   NNPr'  N�r'  h h(h
c__builtin__
__main__
hNN}r'  Ntr'  Rr '  �r!'  Rr"'  NG?�      sX   VBNr#'  ji  �r$'  h h(h
c__builtin__
__main__
hNN}r%'  Ntr&'  Rr''  �r('  Rr)'  (X   TOr*'  G?�=;G ��X   WRBr+'  G?oDe�JBqh�G?�=�	��X   INr,'  G?߬���OX   RBr-'  G?�����i�X   DTr.'  G?��C��,LX   NNr/'  G?��C��,LX   CCr0'  G?�=;G ��X   WPr1'  G?��C��,LX   ''r2'  G?d�C��,LX   JJSr3'  G?d�C��,LX   JJr4'  G?�%����X   RPr5'  G?��C��,LhMG?oDe�JBqX   VBZr6'  G?d�C��,LX   oovr7'  G?d�C��,LX   NNSr8'  G?�=;G ��X   VBGr9'  G?De�JBqX   VBNr:'  G?zT��7^NG?oDe�JBqX   VBPr;'  G?oDe�JBqX   NNPr<'  G?t�C��,LX   ``r='  G?d�C��,Luj
  j�!  �r>'  h h(h
c__builtin__
__main__
hNN}r?'  Ntr@'  RrA'  �rB'  RrC'  (X   VBrD'  G?���B��$h�G?��9��gX   DTrE'  G?��i|Ȯ�X   NNSrF'  G?�K�Ew�`X   NNPrG'  G?���\���X   WPrH'  G?��9��gX   WRBrI'  G?~��Ռ8�X   JJrJ'  G?�K�Ew�`X   PRPrK'  G?���\���X   CDrL'  G?��9��gX   PRP$rM'  G?~��Ռ8�X   RBrN'  G?���\���X   NNrO'  G?���Ռ8�X   VBGrP'  G?���\���X   INrQ'  G?t�9��gX   NNPSrR'  G?t�9��gX   VBNrS'  G?t�9��guj�  j�  �rT'  h h(h
c__builtin__
__main__
hNN}rU'  NtrV'  RrW'  �rX'  RrY'  (X   JJrZ'  G?��l�lX   INr['  G?�`�aX   NNSr\'  G?�X   CCr]'  G?��l�lX   TOr^'  G?�������X   RBr_'  G?�X   NNPr`'  G?��l�lh�G?��l�lX   VBra'  G?��l�lX   NNrb'  G?�X   oovrc'  G?��l�lX   VBGrd'  G?��l�lX   VBNre'  G?�uj\  j  �rf'  h h(h
c__builtin__
__main__
hNN}rg'  Ntrh'  Rri'  �rj'  Rrk'  (h�G?�9GNQӔX   INrl'  G?�
�B�P�X   VBZrm'  G?���+@X   NNrn'  G?�]�a�X   NNPro'  G?�d��!�HX   VBNrp'  G?���+@X   NNSrq'  G?�]�a�X   TOrr'  G?��D��=�X   VBPrs'  G?���+@X   CCrt'  G?�a�AvX   oovru'  G?���+@X   POSrv'  G?���+@X   RBrw'  G?���+@X   VBDrx'  G?���+@X   VBry'  G?����X   JJrz'  G?���+@X   DTr{'  G?����NG?���+@X   ``r|'  G?���+@X   CDr}'  G?����X   WPr~'  G?���+@uX   PRPr'  j�  �r�'  h h(h
c__builtin__
__main__
hNN}r�'  Ntr�'  Rr�'  �r�'  Rr�'  (X   NNPr�'  G?ə�����h�G?�I$�I$�X   POSr�'  G?�A�A�X   CCr�'  G?�A�A�X   ''r�'  G?��_�_X   INr�'  G?�I$�I$�X   VBDr�'  G?�A�A�X   NNr�'  G?�A�A�X   TOr�'  G?��_�_uX   VBNr�'  jj  �r�'  h h(h
c__builtin__
__main__
hNN}r�'  Ntr�'  Rr�'  �r�'  Rr�'  (X   NNSr�'  G?��8�9X   INr�'  G?�-��-��X   TOr�'  G?�W:��th�G?����Q�nX   RBr�'  G?��l�lX   NNr�'  G?�����/X   CCr�'  G?�W:��hMG?�����/hX   VBGr�'  G?�����/hX   JJr�'  G?�q�q�X   NNPr�'  G?�W:��tX   VBPr�'  G?v�l�lX   WRBr�'  G?��l�lX   VBNr�'  G?~W:��tX   WPr�'  G?v�l�lX   ''r�'  G?nW:��tX   WDTr�'  G?nW:��tX   DTr�'  G?nW:��tNG?nW:��tX   VBDr�'  G?nW:��tX   VBr�'  G?nW:��tuhMj�  �r�'  h h(h
c__builtin__
__main__
hNN}r�'  Ntr�'  Rr�'  �r�'  Rr�'  (X   INr�'  G?����i��X   CCr�'  G?���Ez�X   NNPr�'  G?�0ѐX   VBDr�'  G?�2a� &X   MDr�'  G?�0ѐX   RBr�'  G?�0ѐhMG?����i�X   WDTr�'  G?�0ѐX   VBPr�'  G?�0ѐX   TOr�'  G?�0ѐX   NNr�'  G?�0ѐuX   VBNr�'  j�  �r�'  h h(h
c__builtin__
__main__
hNN}r�'  Ntr�'  Rr�'  �r�'  Rr�'  (X   WPr�'  G?�'�n�i�X   NNPr�'  G?����X   INr�'  G?��~�/�RX   TOr�'  G?�n�i�'�h�G?�dI囶X   VBNr�'  G?�yf톙X   PRP$r�'  G?�dI囶X   WRBr�'  G?����Tt X   DTr�'  G?�dI囶X   RBr�'  G?�dI囶X   NNSr�'  G?����Tt X   JJr�'  G?����X   NNr�'  G?����X   JJSr�'  G?����X   CDr�'  G?����X   CCr�'  G?����X   ``r�'  G?����X   oovr�'  G?����Tt X   PRPr�'  G?����Tt X   VBGr�'  G?����uX   WRBr�'  j�  �r�'  h h(h
c__builtin__
__main__
hNN}r�'  Ntr�'  Rr�'  �r�'  Rr�'  (X   VBZr�'  G?خ~G,�tX   NNPr�'  G?�^"p���X   NNSr�'  G?�������X   VBDr�'  G?�����X   INr�'  G?������h�G?������X   RBr�'  G?�^"p���X   MDr�'  G?�^"p���X   NNr�'  G?�8@Ix��X   VBGr�'  G?�^"p���X   CDr�'  G?�^"p���X   CCr�'  G?�^"p���X   VBPr�'  G?��3���jX   JJr�'  G?�^"p���X   NNPSr�'  G?�^"p���X   POSr�'  G?��3���juX   VBDr�'  h_�r�'  h h(h
c__builtin__
__main__
hNN}r�'  Ntr�'  Rr�'  �r�'  Rr�'  (X   NNr�'  G?�}O.��X   NNSr�'  G?�8�13�X   DTr�'  G?�_S˹E�X   VBr�'  G?���;1�PX   NNPr�'  G?�鴩!X   JJr�'  G?������X   INr�'  G?��13��X   RBr�'  G?�sP��'5X   ``r�'  G?x�����X   CDr�'  G?x�����X   PRP$r�'  G?�sP��'5X   VBGr�'  G?����AXiX   WPr�'  G?������h�G?������X   WRBr�'  G?x�����X   POSr�'  G?x�����X   NNPSr�'  G?x�����X   TOr�'  G?��13��hMG?x�����X   RPr�'  G?�sP��'5uX   TOr (  j  �r(  h h(h
c__builtin__
__main__
hNN}r(  Ntr(  Rr(  �r(  Rr(  (X   INr(  G?����hMG?�Y�a�D�h�G?՛�dI�X   RBr(  G?����X   WPr	(  G?����X   PRPr
(  G?u���X   DTr(  G?u���X   VBr(  G?�dI囶X   NNSr(  G?�dI囶X   CCr(  G?����Tt X   VBPr(  G?����Tt X   VBGr(  G?�yf톙X   VBZr(  G?����X   VBDr(  G?����X   TOr(  G?����?WX   VBNr(  G?����Tt X   WDTr(  G?����?WX   NNr(  G?u���X   JJr(  G?u���X   RPr(  G?u���X   NNPr(  G?u���X   WRBr(  G?u���uX   VBZr(  jK  �r(  h h(h
c__builtin__
__main__
hNN}r(  Ntr(  Rr(  �r (  Rr!(  (X   NNr"(  G?�YMe5��X   VBr#(  G?޲��k)�X   JJr$(  G?��SYMe6h�G?�_A}�X   PRPr%(  G?��Gq�wX   NNPr&(  G?��Gq�wX   WPr'(  G?��Gq�wX   NNSr((  G?��w�GqX   TOr)(  G?��_A}�X   INr*(  G?��k)���X   CDr+(  G?��w�GqX   RBr,(  G?��Gq�wX   DTr-(  G?��SYMe6X   CCr.(  G?��w�GqX   VBGr/(  G?��Gq�wX   VBNr0(  G?��Gq�wX   RBSr1(  G?w�_A}�X   PRP$r2(  G?��w�GqX   WRBr3(  G?w�_A}�X   POSr4(  G?w�_A}�X   JJRr5(  G?��Gq�wX   JJSr6(  G?w�_A}�uX   TOr7(  j�  �r8(  h h(h
c__builtin__
__main__
hNN}r9(  Ntr:(  Rr;(  �r<(  Rr=(  (X   VBr>(  G?��;��#�X   INr?(  G?��w�Gqh�G?��SYMe6X   RBr@(  G?��Gq�wX   NNrA(  G?��Gq�wX   CDrB(  G?��Gq�wX   DTrC(  G?��_A}�X   JJrD(  G?��_A}�X   WDTrE(  G?��_A}�X   WPrF(  G?��_A}�hMG?��_A}�X   WRBrG(  G?��_A}�X   VBGrH(  G?��_A}�uX   PRP$rI(  j�  �rJ(  h h(h
c__builtin__
__main__
hNN}rK(  NtrL(  RrM(  �rN(  RrO(  (X   INrP(  G?�I$�I$�X   ''rQ(  G?�I$�I$�X   VBrR(  G?�m��m��X   VBNrS(  G?�m��m��X   JJrT(  G?�I$�I$�ujC  j�  �rU(  h h(h
c__builtin__
__main__
hNN}rV(  NtrW(  RrX(  �rY(  RrZ(  (h�G?��z�-X   INr[(  G?ʧ����lX   TOr\(  G?�+��s��X   JJr](  G?�(��~X   CCr^(  G?�� ��"X   NNr_(  G?�(��~X   MDr`(  G?�$6Qz7X   WPra(  G?�-C���X   VBPrb(  G?�':�Df�X   PRPrc(  G?p$6Qz7X   VBGrd(  G?�*?_��X   VBDre(  G?�(��~X   NNPrf(  G?�$6Qz7X   POSrg(  G?p$6Qz7hMG?�$6Qz7SX   RBrh(  G?�':�Df�X   VBZri(  G?�-C���X   VBNrj(  G?�$6Qz7SX   VBrk(  G?�(��~X   NNSrl(  G?�$6Qz7X   oovrm(  G?�$6Qz7SX   WDTrn(  G?�$6Qz7NG?x$6Qz7SX   DTro(  G?p$6Qz7X   WRBrp(  G?p$6Qz7X   RBSrq(  G?x$6Qz7SuX   INrr(  j8  �rs(  h h(h
c__builtin__
__main__
hNN}rt(  Ntru(  Rrv(  �rw(  Rrx(  (X   RBry(  G?�.)��GXX   PRP$rz(  G?��ͣ��X   VBNr{(  G?�.)��GXX   DTr|(  G?��ͣ��X   CDr}(  G?�.)��GXX   INr~(  G?��ͣ��X   NNPr(  G?��ͣ�X   PRPr�(  G?��y�u�X   WRBr�(  G?�.)��GXX   NNr�(  G?��ͣ�X   VBr�(  G?�.)��GXX   NNSr�(  G?��y�u�X   JJr�(  G?��qO��;X   VBGr�(  G?��qO��;X   TOr�(  G?��qO��;X   ``r�(  G?��qO��;X   JJSr�(  G?��qO��;uj]  j�  �r�(  h h(h
c__builtin__
__main__
hNN}r�(  Ntr�(  Rr�(  �r�(  Rr�(  (X   DTr�(  G?�Y��pȁX   NNPr�(  G?�E�t]FX   VBGr�(  G?�{�D)-X   NNr�(  G?���_X   WPr�(  G?�{�D)-X   JJr�(  G?��;�;X   JJRr�(  G?���^�h�G?���_X   ''r�(  G?�{�D)-X   PRP$r�(  G?�{�D)-X   NNSr�(  G?���_X   INr�(  G?�{�D)-X   PRPr�(  G?���_X   CDr�(  G?���^�X   WRBr�(  G?���^�X   RBr�(  G?�{�D)-X   VBDr�(  G?���^�X   JJSr�(  G?�{�D)-X   WDTr�(  G?�{�D)-X   ``r�(  G?���^�uX   NNPSr�(  h��r�(  h h(h
c__builtin__
__main__
hNN}r�(  Ntr�(  Rr�(  �r�(  Rr�(  (NG?��%VL,X   ``r�(  G?n�ੳӥuX   DTr�(  j�  �r�(  h h(h
c__builtin__
__main__
hNN}r�(  Ntr�(  Rr�(  �r�(  Rr�(  (X   DTr�(  G?��4�,#OX   NNPr�(  G?�i�XF��X   PRP$r�(  G?�{���X   NNSr�(  G?�{���aX   CDr�(  G?��i�XGX   NNr�(  G?��4�,#OX   WDTr�(  G?���a|X   PRPr�(  G?���a|X   JJr�(  G?�a{��X   WPr�(  G?�F��i�X   JJSr�(  G?z{���aX   CCr�(  G?q��a{�X   VBPr�(  G?q��a{�X   JJRr�(  G?q��a{�h�G?���a{�X   INr�(  G?z{���aX   VBGr�(  G?z{���auj  j�  �r�(  h h(h
c__builtin__
__main__
hNN}r�(  Ntr�(  Rr�(  �r�(  Rr�(  (X   INr�(  G?�)ìx�X   JJr�(  G?�~�Q�\X   VBDr�(  G?��� {�	X   VBNr�(  G?ŧ԰V�SX   NNSr�(  G?��԰V�Sh�G?��޾B�{X   VBZr�(  G?���lG'rX   NNr�(  G?��΀b�:X   VBr�(  G?�"ͺd�7X   oovr�(  G?h�΀b�:X   DTr�(  G?���DxX   WPr�(  G?��΀b�:X   VBGr�(  G?���DxX   RBr�(  G?��԰V�SX   MDr�(  G?��԰V�SX   WRBr�(  G?h�΀b�:X   VBPr�(  G?���Po_!X   TOr�(  G?���<S�YX   NNPr�(  G?��԰V�ShMG?��԰V�SX   CCr�(  G?~�� {�	X   ''r�(  G?h�΀b�:X   NNPSr�(  G?h�΀b�:X   PRP$r�(  G?h�΀b�:X   JJSr�(  G?h�΀b�:X   JJRr�(  G?r���J?lX   PRPr�(  G?h�΀b�:uX   WDTr�(  j�  �r�(  h h(h
c__builtin__
__main__
hNN}r�(  Ntr�(  Rr�(  �r�(  Rr�(  (X   VBNr�(  G?�`RjНX   VBDr�(  G?����}�X   NNr�(  G?��|#�9X   NNSr�(  G?������X   RPr�(  G?��n��`RX   INr�(  G?�L��EX   DTr�(  G?Ţ@�´HX   JJr�(  G?��(�0�X   PRPr�(  G?���>X   VBr�(  G?����'%�X   WPr�(  G?��YTy�X   RBr�(  G?�-�Ҭ
MX   JJRr�(  G?��V��X   PRP$r�(  G?��n��`RX   RBSr�(  G?p{�)���X   VBGr�(  G?���>X   TOr�(  G?������X   WRBr�(  G?�{�)���X   NNPr�(  G?��n��`RX   VBZr�(  G?��n��`RX   POSr�(  G?�{�)���h�G?x�n��`RX   VBPr�(  G?p{�)���X   oovr�(  G?x�n��`RX   CCr�(  G?x�n��`RuX   PRP$r )  j�  �r)  h h(h
c__builtin__
__main__
hNN}r)  Ntr)  Rr)  �r)  Rr)  (X   NNr)  G?�+�+�X   JJr)  G?�A�A�X   INr	)  G?�I$�I$�X   RBr
)  G?��_�_X   NNSr)  G?�������h�G?�I$�I$�X   WRBr)  G?�A�A�X   CCr)  G?�A�A�uNh*�r)  h h(h
c__builtin__
__main__
hNN}r)  Ntr)  Rr)  �r)  Rr)  (X   NNr)  G?����E�X   INr)  G?�l2;��qX   TOr)  G?��'��6X   NNSr)  G?�c�{��X   VBDr)  G?�R�+x�X   VBNr)  G?�/U�4*�X   DTr)  G?����[�
hMG?n���E�X   JJr)  G?���<�BX   NNPr)  G?��+x�5"X   POSr)  G?w/U�4*�X   CCr)  G?���<�BX   WPr)  G?���<�BX   MDr )  G?n���E�X   CDr!)  G?w/U�4*�X   VBZr")  G?w/U�4*�X   RBr#)  G?n���E�X   WDTr$)  G?n���E�X   WRBr%)  G?n���E�X   VBGr&)  G?n���E�X   JJRr')  G?n���E�uj|   j�  �r()  h h(h
c__builtin__
__main__
hNN}r))  Ntr*)  Rr+)  �r,)  Rr-)  (X   INr.)  G?���A�JX   VBr/)  G?�X�~��zX   NNr0)  G?�F�eb��X   RBr1)  G?�F�eb��X   VBNr2)  G?�X�~��zX   VBZr3)  G?�F�eb��X   DTr4)  G?��X�~�X   JJr5)  G?�F�eb��X   VBDr6)  G?�F�eb��X   WRBr7)  G?�F�eb��X   NNSr8)  G?�jt�F�X   WDTr9)  G?�F�eb��X   oovr:)  G?�jt�F�uX   DTr;)  j/  �r<)  h h(h
c__builtin__
__main__
hNN}r=)  Ntr>)  Rr?)  �r@)  RrA)  (X   JJrB)  G?ܙɜ�ɝX   VBNrC)  G?���X   RBrD)  G?��J�JX   VBGrE)  G?�A�A�X   NNrF)  G?��Y�YX   JJRrG)  G?���X   CDrH)  G?��h�hX   oovrI)  G?��h�hX   DTrJ)  G?��,�,X   NNSrK)  G?��h�hX   VBPrL)  G?~��X   VBDrM)  G?���X   INrN)  G?~��h�G?��h�hX   TOrO)  G?~��X   VBrP)  G?��,�,X   VBZrQ)  G?��h�hX   NNPrR)  G?~��X   CCrS)  G?~��uNh+�rT)  h h(h
c__builtin__
__main__
hNN}rU)  NtrV)  RrW)  �rX)  RrY)  (X   VBDrZ)  G?���!�xX   NNSr[)  G?�4܁�M�X   VBNr\)  G?�4܁�M�X   INr])  G?�呿YX   VBZr^)  G?�/�A��4X   WDTr_)  G?�% �RPX   VBPr`)  G?�4܁�M�X   MDra)  G?�4܁�M�X   NNPrb)  G?~4܁�M�X   VBGrc)  G?���ajzVX   RBrd)  G?�*J���X   CCre)  G?���ajzVX   WPrf)  G?����X   TOrg)  G?����X   JJrh)  G?���	�.X   oovri)  G?h*J���hMG?���!�xX   POSrj)  G?x*J���X   VBrk)  G?~4܁�M�X   RBSrl)  G?h*J���X   JJRrm)  G?h*J���X   DTrn)  G?r��!�xX   NNro)  G?~4܁�M�X   WRBrp)  G?h*J���uX   CDrq)  j�
  �rr)  h h(h
c__builtin__
__main__
hNN}rs)  Ntrt)  Rru)  �rv)  Rrw)  (X   NNSrx)  G?�333333h�G?�333333hMG?�������X   JJry)  G?�������X   WPrz)  G?�333333X   NNr{)  G?�      X   CCr|)  G?�������X   INr})  G?�333333X   NNPr~)  G?�������X   VBDr)  G?�      X   JJRr�)  G?�333333X   WRBr�)  G?�������X   PRPr�)  G?�������X   TOr�)  G?�������X   NNPSr�)  G?�������X   VBNr�)  G?�������X   DTr�)  G?�������uX   PRPr�)  j�  �r�)  h h(h
c__builtin__
__main__
hNN}r�)  Ntr�)  Rr�)  �r�)  Rr�)  (X   VBr�)  G?�������X   NNPr�)  G?�ffffffh�G?�������X   WPr�)  G?�      X   DTr�)  G?�ffffffX   PRPr�)  G?�������X   RBr�)  G?�������X   JJr�)  G?�������X   NNSr�)  G?�������X   INr�)  G?�333333X   ``r�)  G?�������X   CDr�)  G?�������uX   VBPr�)  j�  �r�)  h h(h
c__builtin__
__main__
hNN}r�)  Ntr�)  Rr�)  �r�)  Rr�)  (X   NNSr�)  G?������X   INr�)  G?ы�YR$�hMG?�z��q?X   VBGr�)  G?���YR$�X   NNr�)  G?��C���h�G?ƺ��#�X   CCr�)  G?��/���X   TOr�)  G?���"J�X   WRBr�)  G?y�/���X   VBDr�)  G?�T�+���X   MDr�)  G?y�/���X   VBZr�)  G?��/���X   JJRr�)  G?i�/���X   VBPr�)  G?s#�J+�X   VBNr�)  G?����@�X   WDTr�)  G?y�/���X   ''r�)  G?y�/���X   PRPr�)  G?s#�J+�X   RBr�)  G?�T�+���X   VBr�)  G?y�/���X   POSr�)  G?�T�+���X   JJr�)  G?y�/���X   DTr�)  G?i�/���X   NNPr�)  G?i�/���NG?i�/���X   WPr�)  G?s#�J+�X   CDr�)  G?i�/���uj1	  hM�r�)  h h(h
c__builtin__
__main__
hNN}r�)  Ntr�)  Rr�)  �r�)  Rr�)  (X   NNPr�)  G?��o��o�X   WRBr�)  G?� � �X   VBGr�)  G?�A�A�X   VBZr�)  G?��;�;X   WDTr�)  G?��;�;X   NNSr�)  G?�A�A�X   WPr�)  G?�-��-��X   INr�)  G?�A�A�X   JJr�)  G?�A�A�X   NNr�)  G?��;�;X   ''r�)  G?��;�;X   DTr�)  G?��؝�؞X   PRPr�)  G?�i�i�X   VBr�)  G?�A�A�X   VBNr�)  G?�A�A�X   MDr�)  G?��;�;X   CCr�)  G?��؝�؞X   VBDr�)  G?�A�A�X   RBr�)  G?�i�i�X   VBPr�)  G?��;�;X   CDr�)  G?�A�A�ujl  jV  �r�)  h h(h
c__builtin__
__main__
hNN}r�)  Ntr�)  Rr�)  �r�)  Rr�)  (X   NNPr�)  G?�i�i�X   WPr�)  G?�A�A�X   DTr�)  G?��;�;X   CDr�)  G?� � �X   JJr�)  G?�A�A�X   POSr�)  G?�A�A�X   NNr�)  G?�A�A�X   VBZr�)  G?�A�A�X   PRP$r�)  G?��;�;uX   CCr�)  j�  �r�)  h h(h
c__builtin__
__main__
hNN}r�)  Ntr�)  Rr�)  �r�)  Rr�)  (X   VBDr�)  G?�?����X   VBPr�)  G?�h�G?ӷy;phX   INr�)  G?��J���X   NNr�)  G?�\��eϾX   VBZr�)  G?���!�y�X   TOr�)  G?�ǀ��xX   VBNr�)  G?��L�x��X   JJr�)  G?���a{�hMG?��7Q�cuX   oovr�)  G?w�L�x��X   NNPr�)  G?b�
-P�X   RBr�)  G?�\��eϾX   CCr�)  G?�zh���X   VBr�)  G?�/�AR��X   JJRr�)  G?l?����X   VBGr�)  G?|?����X   MDr�)  G?|?����X   WDTr�)  G?��L�x��X   RBSr�)  G?r�
-P�X   DTr�)  G?|?����X   POSr�)  G?l?����X   WPr�)  G?l?����X   ''r�)  G?l?����X   NNSr�)  G?�/�AR��X   CDr *  G?b�
-P�X   PRPr*  G?b�
-P�NG?l?����X   RPr*  G?b�
-P�uX   MDr*  j"  �r*  h h(h
c__builtin__
__main__
hNN}r*  Ntr*  Rr*  �r*  Rr	*  (X   JJr
*  G?�Ӹ�<X   NNr*  G?�����YX   NNPr*  G?Ë�8�X   NNSr*  G?�L���X   JJRr*  G?�_{(!5�X   VBGr*  G?�#�wb@X   CDr*  G?��y�ᎈX   INr*  G?����A	�X   VBr*  G?�_{(!5�X   VBNr*  G?�#�wb@X   oovr*  G?v#�wb@X   ``r*  G?p���A	�X   RBr*  G?��y�ᎈX   JJSr*  G?v#�wb@X   NNPSr*  G?f#�wb@X   RBSr*  G?f#�wb@uX   CCr*  j�  �r*  h h(h
c__builtin__
__main__
hNN}r*  Ntr*  Rr*  �r*  Rr *  (X   INr!*  G?�E�t]FX   JJr"*  G?ދ��.�X   VBPr#*  G?�]E�t]X   NNr$*  G?�E�t]FX   NNSr%*  G?�t]E�tX   VBZr&*  G?�t]E�tuj�  j!*  �r'*  h h(h
c__builtin__
__main__
hNN}r(*  Ntr)*  Rr**  �r+*  Rr,*  (X   NNPr-*  G?�;�6w�mX   DTr.*  G?�Ɉ+�X   PRP$r/*  G?�W& �LAX   JJr0*  G?�Ɉ+�WX   CDr1*  G?�Ɉ+�WX   VBGr2*  G?�Ɉ+�WX   JJSr3*  G?�W& �LAuX   NNSr4*  j@  �r5*  h h(h
c__builtin__
__main__
hNN}r6*  Ntr7*  Rr8*  �r9*  Rr:*  (X   PRPr;*  G?��/�A�3X   VBr<*  G?�A�l'TX   RBr=*  G?�8d���X   DTr>*  G?�O�豴�X   NNr?*  G?�8d���X   JJr@*  G?wNKt�X   NNPrA*  G?��/�A�3X   NNSrB*  G?�NKt�X   CDrC*  G?�z�C�X   VBGrD*  G?wNKt�X   VBDrE*  G?qz�C�X   WPrF*  G?wNKt�h�G?wNKt�X   PRP$rG*  G?gNKt�X   INrH*  G?qz�C�X   VBNrI*  G?gNKt�uX   CDrJ*  j�
  �rK*  h h(h
c__builtin__
__main__
hNN}rL*  NtrM*  RrN*  �rO*  RrP*  (X   VBDrQ*  G?斖����X   VBNrR*  G?�X   NNSrS*  G?�X   NNPrT*  G?�������X   NNrU*  G?�������X   VBZrV*  G?�X   VBPrW*  G?�X   JJrX*  G?�X   RBrY*  G?�uj�  j�  �rZ*  h h(h
c__builtin__
__main__
hNN}r[*  Ntr\*  Rr]*  �r^*  Rr_*  (X   VBDr`*  G?���q�X   NNSra*  G?�+���^X   VBZrb*  G?�����X   MDrc*  G?�5���*X   VBPrd*  G?���6��X   NNPre*  G?�v��K,X   CDrf*  G?p��sl�X   NNrg*  G?���jY_�X   RBrh*  G?��`M���X   TOri*  G?f+���^X   JJrj*  G?�v��K,X   WPrk*  G?f+���^X   JJSrl*  G?f+���^X   DTrm*  G?p��sl�X   oovrn*  G?p��sl�X   INro*  G?p��sl�uX   WPrp*  jk  �rq*  h h(h
c__builtin__
__main__
hNN}rr*  Ntrs*  Rrt*  �ru*  Rrv*  (X   VBrw*  G?�1Yr��X   PRPrx*  G?���k�X   DTry*  G?Ȭ�k�X   NNSrz*  G?��!�~u4X   PRP$r{*  G?���k�X   JJr|*  G?���k�X   NNr}*  G?���k�X   NNPr~*  G?���k�uj�  je  �r*  h h(h
c__builtin__
__main__
hNN}r�*  Ntr�*  Rr�*  �r�*  Rr�*  (X   VBDr�*  G?�X   INr�*  G?ϱ��� h�G?ĹK��K�X   RBr�*  G?�A�A�X   WPr�*  G?��8�8X   VBPr�*  G?��_�_X   NNr�*  G?��8�8X   TOr�*  G?��8�8hMG?��8�8X   DTr�*  G?�A�A�X   NNPr�*  G?��8�8X   POSr�*  G?��8�8X   WRBr�*  G?��8�8X   NNSr�*  G?��8�8X   MDr�*  G?�A�A�X   VBr�*  G?��8�8X   VBNr�*  G?��8�8X   NNPSr�*  G?��8�8X   VBGr�*  G?��8�8uX   INr�*  j�  �r�*  h h(h
c__builtin__
__main__
hNN}r�*  Ntr�*  Rr�*  �r�*  Rr�*  (X   VBr�*  G?� �� ��X   NNPr�*  G?�^�^�X   DTr�*  G?�����h�G?��$�$X   CCr�*  G?�����X   RBr�*  G?�~h~hX   WPr�*  G?�~h~hX   PRP$r�*  G?�~h~hX   NNr�*  G?�����X   INr�*  G?�>�>�X   WRBr�*  G?�����X   oovr�*  G?�����X   JJr�*  G?�����X   CDr�*  G?�~h~hX   VBGr�*  G?�~h~hX   WDTr�*  G?�����X   NNSr�*  G?�����uhMj.  �r�*  h h(h
c__builtin__
__main__
hNN}r�*  Ntr�*  Rr�*  �r�*  Rr�*  (X   NNPr�*  G?�#��`�X   JJr�*  G?�#��`�X   NNr�*  G?�a����X   VBNr�*  G?�bM���X   VBZr�*  G?�N���OX   NNSr�*  G?�5�@+��X   JJRr�*  G?�bM���X   INr�*  G?�bM���X   RBSr�*  G?�bM���X   NNPSr�*  G?�Z�oFQX   VBGr�*  G?u�g���X   RBr�*  G?�bM���hMG?�bM���X   CDr�*  G?�bM���X   JJSr�*  G?�bM���X   VBPr�*  G?�bM���uj�  j�  �r�*  h h(h
c__builtin__
__main__
hNN}r�*  Ntr�*  Rr�*  �r�*  Rr�*  (X   INr�*  G?��Z��Eh�G?��� ��TX   TOr�*  G?�=��X�X   VBr�*  G?�R�+x�X   VBPr�*  G?��7ܷ��X   RBr�*  G?��7ܷ��X   WRBr�*  G?j�~�N�X   VBNr�*  G?�@p�X   JJr�*  G?�{�4�JX   VBDr�*  G?��h_Ä�X   NNr�*  G?~=��X�hMG?�{�4�JX   NNSr�*  G?d))_";9X   VBGr�*  G?�=��X�X   VBZr�*  G?�R�+x�X   JJSr�*  G?Z�~�N�X   oovr�*  G?~=��X�X   DTr�*  G?�{�4�JX   NNPr�*  G?j�~�N�X   CCr�*  G?p���G1ZX   PRP$r�*  G?j�~�N�X   MDr�*  G?Z�~�N�X   JJRr�*  G?d))_";9NG?Z�~�N�X   WPr�*  G?Z�~�N�X   RPr�*  G?d))_";9X   CDr�*  G?Z�~�N�X   ``r�*  G?Z�~�N�ujf  j�  �r�*  h h(h
c__builtin__
__main__
hNN}r�*  Ntr�*  Rr�*  �r�*  Rr�*  (X   NNPr�*  G?��~2z�pX   NNSr�*  G?��d�.ߍX   NNr�*  G?��d�.ߍX   JJr�*  G?�z�o�OSX   VBGr�*  G?|�V��X   NNPSr�*  G?|�V��X   CDr�*  G?��@�´Hh�G?|�V��X   JJRr�*  G?�6�@�X   VBDr�*  G?|�V��X   JJSr�*  G?|�V��X   VBNr�*  G?|�V��X   RBr�*  G?��@�´HuX   VBr�*  j*  �r�*  h h(h
c__builtin__
__main__
hNN}r�*  Ntr�*  Rr�*  �r�*  Rr�*  (X   NNPr�*  G?�^rT�>#X   JJr�*  G?�e�%HX   VBDr�*  G?��,��X   DTr�*  G?��CV��X   VBNr�*  G?��CV��X   NNSr�*  G?��,��X   NNr +  G?�^rT�>#X   RBr+  G?�ڷ��CX   PRP$r+  G?��,��X   oovr+  G?��,��h�G?�V���hcX   VBr+  G?�ڷ��CX   CCr+  G?��,��X   CDr+  G?��,��X   MDr+  G?��CV��uX   VBZr+  jL  �r	+  h h(h
c__builtin__
__main__
hNN}r
+  Ntr+  Rr+  �r+  Rr+  (X   TOr+  G?�X��Ƈ�X   VBr+  G?�8N��X   VBNr+  G?�j;5��[h�G?��+���X   DTr+  G?����kdmX   WPr+  G?�AAX   RBr+  G?��r[��X   INr+  G?��5g�ǱX   NNr+  G?�z|:�_X   NNSr+  G?���c؆�X   JJr+  G?�a�a�X   VBDr+  G?r�r[��X   CCr+  G?�8N��X   PRPr+  G?��r[��hMG?��r[��X   POSr+  G?��r[��X   NNPr+  G?����s��X   VBZr+  G?r�r[��X   oovr+  G?��r[��X   JJRr +  G?{�+���X   CDr!+  G?{�+���X   RPr"+  G?�8N��X   PRP$r#+  G?{�+���NG?r�r[��X   VBGr$+  G?{�+���X   ''r%+  G?��r[��X   WRBr&+  G?{�+���uX   CDr'+  jM  �r(+  h h(h
c__builtin__
__main__
hNN}r)+  Ntr*+  Rr++  �r,+  Rr-+  (X   VBDr.+  G?˻�����X   JJr/+  G?�X   RBr0+  G?�������X   NNPr1+  G?�X   PRPr2+  G?�X   DTr3+  G?�������X   NNr4+  G?�uj�   j3#  �r5+  h h(h
c__builtin__
__main__
hNN}r6+  Ntr7+  Rr8+  �r9+  Rr:+  (X   PRPr;+  G?�;�;�X   VBGr<+  G?��؝�؞X   VBNr=+  G?��;�;X   NNSr>+  G?ȝ�؝��X   DTr?+  G?ñ;�;X   VBDr@+  G?��؝�؞X   NNrA+  G?��;�;uh�j�  �rB+  h h(h
c__builtin__
__main__
hNN}rC+  NtrD+  RrE+  �rF+  RrG+  (h�G?ݶ�m��nX   NNPrH+  G?�I$�I$�hMG?�I$�I$�NG?�m��m��X   INrI+  G?�I$�I$�uj�  h��rJ+  h h(h
c__builtin__
__main__
hNN}rK+  NtrL+  RrM+  �rN+  RrO+  NG?�      sX   WPrP+  j  �rQ+  h h(h
c__builtin__
__main__
hNN}rR+  NtrS+  RrT+  �rU+  RrV+  (X   NNrW+  G?�UUUUUUX   TOrX+  G?�      X   VBDrY+  G?��8�9X   VBNrZ+  G?�q�q�X   JJr[+  G?��8�9X   POSr\+  G?�q�q�X   NNSr]+  G?�q�q�X   VBGr^+  G?�q�q�X   INr_+  G?��8�9X   RPr`+  G?�q�q�X   DTra+  G?�q�q�X   VBZrb+  G?�q�q�X   NNPrc+  G?�UUUUUUX   RBrd+  G?�q�q�X   MDre+  G?�q�q�X   VBPrf+  G?�q�q�uX   VBGrg+  j�	  �rh+  h h(h
c__builtin__
__main__
hNN}ri+  Ntrj+  Rrk+  �rl+  Rrm+  (X   DTrn+  G?͉؝�؞X   WDTro+  G?�A�A�X   NNPrp+  G?� � �X   VBNrq+  G?�A�A�X   NNrr+  G?�A�A�X   RBrs+  G?�i�i�X   INrt+  G?��o��o�X   TOru+  G?��o��o�X   JJrv+  G?�A�A�X   WPrw+  G?�A�A�X   PRPrx+  G?�A�A�X   CCry+  G?��;�;X   RPrz+  G?�A�A�h�G?�A�A�X   JJRr{+  G?�A�A�X   NNSr|+  G?��;�;uX   CCr}+  j�  �r~+  h h(h
c__builtin__
__main__
hNN}r+  Ntr�+  Rr�+  �r�+  Rr�+  (h�G?̕ O���X   PRPr�+  G?��,��X   INr�+  G?�^rT�>#hMG?��CV��X   TOr�+  G?�ڷ��CX   JJr�+  G?�ڷ��CX   NNSr�+  G?�e�%H�X   NNr�+  G?�'�Yy�RX   CCr�+  G?��CV��X   DTr�+  G?�ڷ��CX   WRBr�+  G?��,��X   RBr�+  G?��,��X   NNPr�+  G?��CV��X   VBGr�+  G?��,��X   WPr�+  G?��CV��X   RPr�+  G?��,��X   JJRr�+  G?��CV��X   oovr�+  G?��,��X   VBNr�+  G?��,��uj�  j  �r�+  h h(h
c__builtin__
__main__
hNN}r�+  Ntr�+  Rr�+  �r�+  Rr�+  (X   WRBr�+  G?��a���X   RPr�+  G?��A)��X   INr�+  G?A)��X   NNPr�+  G?��A)��X   VBGr�+  G?��A)��X   VBNr�+  G?��A)��X   NNSr�+  G?�E�t]FX   DTr�+  G?�Jy��Jh�G?��A)��X   JJr�+  G?��A)��X   JJSr�+  G?��A)��X   CCr�+  G?��A)��X   TOr�+  G?��A)��hMG?��A)��X   WPr�+  G?��A)��X   NNr�+  G?��A)��uj  j�+  �r�+  h h(h
c__builtin__
__main__
hNN}r�+  Ntr�+  Rr�+  �r�+  Rr�+  (X   PRPr�+  G?Ҍ�J3�)X   RBr�+  G?��`v���h�G?�B�Y!dX   JJr�+  G?�J3�)X   DTr�+  G?��B�YX   NNPr�+  G?�B�Y!dX   NNr�+  G?��`v���X   TOr�+  G?�B�Y!dX   VBNr�+  G?�B�Y!dX   VBDr�+  G?��`v���X   VBGr�+  G?���J3�)X   NNSr�+  G?��`v���X   oovr�+  G?��`v���uX   NNSr�+  jA  �r�+  h h(h
c__builtin__
__main__
hNN}r�+  Ntr�+  Rr�+  �r�+  Rr�+  (X   VBDr�+  G?�333333X   VBPr�+  G?��_�_X   DTr�+  G?�A�A�X   MDr�+  G?�uPuPX   VBZr�+  G?�I$�I$�X   RBr�+  G?��_�_X   INr�+  G?�uPuPX   TOr�+  G?�A�A�X   VBGr�+  G?�A�A�uX   NNr�+  j3	  �r�+  h h(h
c__builtin__
__main__
hNN}r�+  Ntr�+  Rr�+  �r�+  Rr�+  (X   VBDr�+  G?����{��X   NNPr�+  G?�D�4MEX   VBZr�+  G?�7�p�7X   NNr�+  G?�4MD�4X   RBr�+  G?�e�v]�fh�G?���n�X   PRPr�+  G?��!B�X   MDr�+  G?��9�s��X   JJr�+  G?���n�X   VBPr�+  G?���n�X   INr�+  G?��`XhMG?v�`XX   WRBr�+  G?v�`XX   CDr�+  G?v�`XX   NNSr�+  G?v�`Xuj�  jZ  �r�+  h h(h
c__builtin__
__main__
hNN}r�+  Ntr�+  Rr�+  �r�+  Rr�+  X   RBr�+  G?�      sX   VBPr�+  jJ  �r�+  h h(h
c__builtin__
__main__
hNN}r�+  Ntr�+  Rr�+  �r�+  Rr�+  (X   NNSr�+  G?�b�b�b�X   JJr�+  G?����X   TOr�+  G?���� X   INr�+  G?����X   RBr�+  G?��� X   NNr�+  G?����X   CCr�+  G?����X   JJRr�+  G?��� h�G?���� X   NNPr�+  G?���� X   DTr�+  G?��� X   VBGr�+  G?��� X   CDr�+  G?����hMG?��� ujC)  j+  �r�+  h h(h
c__builtin__
__main__
hNN}r�+  Ntr�+  Rr�+  �r�+  Rr�+  (h�G?�����/hX   RBr�+  G?�q�q�X   DTr ,  G?�����/hX   INr,  G?���%�	{X   JJr,  G?�����/huj+  h��r,  h h(h
c__builtin__
__main__
hNN}r,  Ntr,  Rr,  �r,  Rr,  NG?�      sX   VBNr	,  j�  �r
,  h h(h
c__builtin__
__main__
hNN}r,  Ntr,  Rr,  �r,  Rr,  (X   NNr,  G?��� U9X   JJr,  G?Πu.E�X   NNPr,  G?��T9B?X   JJSr,  G?����h3X   WPr,  G?�N;A��fX   RBSr,  G?��X7�[�X   VBGr,  G?�N;A��fX   NNSr,  G?���U�&X   VBNr,  G?eN;A��fX   ``r,  G?��s�b4�X   oovr,  G?uN;A��fX   DTr,  G?�N;A��fX   INr,  G?�����X   CDr,  G?�X�_5�X   VBZr,  G?��s�b4�X   JJRr,  G?uN;A��fX   RBr ,  G?uN;A��fX   MDr!,  G?uN;A��fX   VBPr",  G?eN;A��fX   VBDr#,  G?eN;A��fX   VBr$,  G?eN;A��fNG?eN;A��fuX   VBr%,  h��r&,  h h(h
c__builtin__
__main__
hNN}r',  Ntr(,  Rr),  �r*,  Rr+,  (X   INr,,  G?�Pה5�X   NNSr-,  G?ǔ5�yCX   NNr.,  G?�򆼡�(X   JJr/,  G?�򆼡�(X   RBr0,  G?�򆼡�(X   TOr1,  G?�򆼡�(h�G?�5�yC^uX   POSr2,  jW  �r3,  h h(h
c__builtin__
__main__
hNN}r4,  Ntr5,  Rr6,  �r7,  Rr8,  (X   NNSr9,  G?�
�cp"X   NNr:,  G?ˁ�V�jX   INr;,  G?�7��}X   JJr<,  G?�cp!���X   TOr=,  G?�(2��C�X   WPr>,  G?���k朐h�G?ӑ��¥X   VBZr?,  G?���k朐X   RPr@,  G?�cp!���X   CCrA,  G?���k朐X   NNPrB,  G?���k朐X   VBPrC,  G?���k朐X   VBDrD,  G?���k朐X   VBNrE,  G?���k朐uX   VBPrF,  j
  �rG,  h h(h
c__builtin__
__main__
hNN}rH,  NtrI,  RrJ,  �rK,  RrL,  (h�G?�~��TxX   NNrM,  G?٪;�҄�X   RBrN,  G?�ʸ�%�nX   NNPrO,  G?�0ʸ�&X   TOrP,  G?�d�
e\X   CDrQ,  G?�ʸ�%�nX   INrR,  G?������8X   oovrS,  G?�ʸ�%�nX   VBZrT,  G?�ʸ�%�nX   JJrU,  G?�d�
e\X   NNSrV,  G?��f��JX   MDrW,  G?�ʸ�%�nX   DTrX,  G?�ʸ�%�nuhMj�  �rY,  h h(h
c__builtin__
__main__
hNN}rZ,  Ntr[,  Rr\,  �r],  Rr^,  (X   INr_,  G?�X   NNr`,  G?�������X   NNSra,  G?�ffffffhMG?�""""""h�G?�������X   CCrb,  G?�DDDDDDX   ``rc,  G?�X   VBZrd,  G?�wwwwwwX   TOre,  G?�UUUUUUX   RBrf,  G?y������X   ''rg,  G?y������X   NNPrh,  G?�X   MDri,  G?�������X   VBDrj,  G?�������X   CDrk,  G?�X   VBNrl,  G?qX   JJrm,  G?qX   PRPrn,  G?qX   DTro,  G?y������X   VBGrp,  G?qX   JJRrq,  G?quj�  j�%  �rr,  h h(h
c__builtin__
__main__
hNN}rs,  Ntrt,  Rru,  �rv,  Rrw,  (X   INrx,  G?�<<<<<<X   NNSry,  G?�������h�G?д�����X   VBZrz,  G?�������X   TOr{,  G?�������X   NNr|,  G?�<<<<<<X   VBr},  G?�X   WDTr~,  G?~X   WPr,  G?�X   CCr�,  G?�X   VBNr�,  G?�������X   RBr�,  G?�������X   JJr�,  G?�X   WRBr�,  G?�������X   VBDr�,  G?�X   DTr�,  G?�X   ''r�,  G?~X   oovr�,  G?~X   MDr�,  G?~X   JJRr�,  G?~hMG?~X   NNPr�,  G?~uX   WRBr�,  j  �r�,  h h(h
c__builtin__
__main__
hNN}r�,  Ntr�,  Rr�,  �r�,  Rr�,  (X   NNr�,  G?�I$�I$�X   NNSr�,  G?�I$�I$�X   VBNr�,  G?�I$�I$�uX   JJSr�,  j  �r�,  h h(h
c__builtin__
__main__
hNN}r�,  Ntr�,  Rr�,  �r�,  Rr�,  (X   JJr�,  G?�+��Q,X   NNr�,  G?�+��Q,X   NNPr�,  G?������X   INr�,  G?������X   NNSr�,  G?������uj
  j�  �r�,  h h(h
c__builtin__
__main__
hNN}r�,  Ntr�,  Rr�,  �r�,  Rr�,  (X   DTr�,  G?�]~��&X   JJr�,  G?�B�Y!dX   RBr�,  G?���s��X   oovr�,  G?�����X   VBGr�,  G?�����X   VBNr�,  G?�����X   JJRr�,  G?�����X   NNr�,  G?�*K��a�X   INr�,  G?���s��X   NNPr�,  G?���s��X   CCr�,  G?�����h�G?���s��X   VBDr�,  G?�����uX   INr�,  hM�r�,  h h(h
c__builtin__
__main__
hNN}r�,  Ntr�,  Rr�,  �r�,  Rr�,  (X   VBNr�,  G?��O��X   CCr�,  G?���`jc�X   NNr�,  G?���`jc�X   RBr�,  G?��O��X   WPr�,  G?��Lw�5X   INr�,  G?՜B~Vq
X   NNSr�,  G?��O��X   WDTr�,  G?���`jc�X   TOr�,  G?���`jc�X   NNPr�,  G?���`jc�X   VBGr�,  G?���`jc�X   PRPr�,  G?���`jc�X   DTr�,  G?���`jc�uX   VBNr�,  j�  �r�,  h h(h
c__builtin__
__main__
hNN}r�,  Ntr�,  Rr�,  �r�,  Rr�,  (X   INr�,  G?ڙϊdhMG?�� ��F�h�G?�� ��GX   TOr�,  G?�y&���X   DTr�,  G?�d�ҳX   WDTr�,  G?�� ��F�X   NNPr�,  G?�� ��F�X   VBGr�,  G?��ҳ;X   WRBr�,  G?�H�����X   RBr�,  G?�H�����X   JJr�,  G?�H�����X   oovr�,  G?�� ��F�X   NNSr�,  G?�� ��F�X   WPr�,  G?�H�����X   NNr�,  G?�H�����X   CDr�,  G?�� ��F�uX   TOr�,  jF!  �r�,  h h(h
c__builtin__
__main__
hNN}r�,  Ntr�,  Rr�,  �r�,  Rr�,  (h�G?̼��/X   VBGr�,  G?�I$�I$�X   JJr�,  G?ѡ���hX   VBDr�,  G?�X��ƈX   NNr�,  G?���/9X   INr�,  G?���/9X   PRPr�,  G?�X��ƈX   DTr�,  G?�X��ƈX   RBr�,  G?���/9X   JJRr�,  G?���/9X   VBZr�,  G?���/9X   VBNr�,  G?�X��Ƈ�X   MDr�,  G?���/9X   VBPr�,  G?���/9uX   NNSr�,  j�  �r�,  h h(h
c__builtin__
__main__
hNN}r�,  Ntr�,  Rr�,  �r�,  Rr�,  (X   VBDr�,  G?����X   NNr�,  G?���^�X   VBPr�,  G?��}P�X   WPr�,  G?|��^�h�G?�E�t]FX   VBZr�,  G?���_X   JJr�,  G?�{�D)-hMG?�{�D)-X   RBr�,  G?����[L�X   MDr�,  G?�{�D)-NG?|��^�X   NNSr -  G?|��^�X   CDr-  G?|��^�X   PRPr-  G?|��^�X   VBr-  G?|��^�X   INr-  G?|��^�X   DTr-  G?|��^�uX   WRBr-  j�  �r-  h h(h
c__builtin__
__main__
hNN}r-  Ntr	-  Rr
-  �r-  Rr-  (X   VBr-  G?�>���>X   NNr-  G?���|X   WRBr-  G?���|X   RBr-  G?���|uX   JJr-  j�  �r-  h h(h
c__builtin__
__main__
hNN}r-  Ntr-  Rr-  �r-  Rr-  (X   JJr-  G?��Ҽy�XX   NNr-  G?�J���a5X   VBNr-  G?ə�����X   INr-  G?�J3�)h�G?��V�AX   RBr-  G?�J���a5X   TOr-  G?�B�Y!dX   VBDr-  G?�*K��a�hMG?��`v���X   VBZr-  G?�*K��a�X   DTr -  G?��`v���X   VBGr!-  G?�����X   VBr"-  G?�����X   NNSr#-  G?����ALX   NNPr$-  G?��`v���X   WRBr%-  G?�����X   ''r&-  G?w���.|X   oovr'-  G?�����X   CCr(-  G?w���.|X   VBPr)-  G?����ALX   MDr*-  G?�����uhMj�  �r+-  h h(h
c__builtin__
__main__
hNN}r,-  Ntr--  Rr.-  �r/-  Rr0-  (X   RPr1-  G?�UUUUUUh�G?�I$�I$�X   NNr2-  G?�y�y�X   TOr3-  G?�I$�I$�X   RBr4-  G?�a�a�X   NNSr5-  G?�I$�I$�X   CCr6-  G?�I$�I$�X   NNPr7-  G?�a�a�hMG?�a�a�X   VBNr8-  G?�a�a�X   PRP$r9-  G?�a�a�X   PRPr:-  G?�a�a�X   WRBr;-  G?�a�a�uNh,�r<-  h h(h
c__builtin__
__main__
hNN}r=-  Ntr>-  Rr?-  �r@-  RrA-  (X   DTrB-  G?�!d,���X   PRPrC-  G?��zoM�X   RBrD-  G?�B�Y!duX   VBNrE-  j   �rF-  h h(h
c__builtin__
__main__
hNN}rG-  NtrH-  RrI-  �rJ-  RrK-  (X   INrL-  G?���5_�X   VBNrM-  G?����X   TOrN-  G?�4b�y�Fh�G?�� �%�RhMG?���J!�.X   JJrO-  G?���/q��X   RBrP-  G?�ʠ��X   PRPrQ-  G?w���{�X   WRBrR-  G?w���{�X   CDrS-  G?w���{�X   NNSrT-  G?o���X   VBGrU-  G?�ʠ��X   DTrV-  G?����{�X   VBrW-  G?����{�X   oovrX-  G?w���{�X   VBZrY-  G?w���{�X   CCrZ-  G?������X   JJRr[-  G?w���{�X   WDTr\-  G?o���X   NNr]-  G?���X   NNPr^-  G?o���X   VBDr_-  G?o���X   PRP$r`-  G?o���uh�j�  �ra-  h h(h
c__builtin__
__main__
hNN}rb-  Ntrc-  Rrd-  �re-  Rrf-  (X   INrg-  G?�      h�G?�I$�I$�X   NNSrh-  G?�I$�I$�hMG?��m��m�X   VBZri-  G?�I$�I$�X   VBNrj-  G?��m��m�X   NNPrk-  G?�I$�I$�X   VBPrl-  G?�I$�I$�X   CCrm-  G?�m��m��X   JJrn-  G?�I$�I$�X   oovro-  G?�I$�I$�NG?�I$�I$�X   VBDrp-  G?�I$�I$�X   NNrq-  G?�m��m��uX   VBrr-  h��rs-  h h(h
c__builtin__
__main__
hNN}rt-  Ntru-  Rrv-  �rw-  Rrx-  (X   PRPry-  G?�UUUUUUX   PRP$rz-  G?�X   RBr{-  G?�X   VBGr|-  G?�������X   JJr}-  G?�PPPPPPX   DTr~-  G?�������X   NNSr-  G?�������h�G?�������X   NNr�-  G?�X   VBNr�-  G?�X   INr�-  G?�������X   VBr�-  G?�X   NNPr�-  G?�X   WPr�-  G?�X   CDr�-  G?�X   TOr�-  G?�X   RPr�-  G?�uX   RPr�-  j�  �r�-  h h(h
c__builtin__
__main__
hNN}r�-  Ntr�-  Rr�-  �r�-  Rr�-  (X   INr�-  G?�UUUUUUh�G?�UUUUUUX   VBDr�-  G?�UUUUUUuj�  j�-  �r�-  h h(h
c__builtin__
__main__
hNN}r�-  Ntr�-  Rr�-  �r�-  Rr�-  (X   DTr�-  G?��	�}�X   JJr�-  G?��`����X   NNr�-  G?�eo&�:X   NNPr�-  G?ć>��0MX   CCr�-  G?�R�+x�X   VBNr�-  G?��+x�5"X   INr�-  G?�&�9�V�X   ''r�-  G?��+x�5"X   ``r�-  G?��`����X   NNSr�-  G?�R�+x�X   oovr�-  G?��+x�5"X   PRP$r�-  G?���[�	�X   PRPr�-  G?��+x�5"uj^  j�  �r�-  h h(h
c__builtin__
__main__
hNN}r�-  Ntr�-  Rr�-  �r�-  Rr�-  (X   VBNr�-  G?�A�A�X   NNSr�-  G?��_�_X   TOr�-  G?��_�_X   INr�-  G?�uPuPX   VBGr�-  G?�A�A�X   NNr�-  G?�I$�I$�X   NNPr�-  G?�A�A�X   JJr�-  G?�������X   NNPSr�-  G?�A�A�h�G?�A�A�uj6	  j�  �r�-  h h(h
c__builtin__
__main__
hNN}r�-  Ntr�-  Rr�-  �r�-  Rr�-  (X   VBGr�-  G?��+���X   PRP$r�-  G?��+���X   NNPr�-  G?�m��m��X   DTr�-  G?���{�qX   NNSr�-  G?�j;5��[X   JJr�-  G?�j;5��[X   VBPr�-  G?��+���X   NNr�-  G?�X��Ƈ�X   CDr�-  G?���/9h�G?��+���X   INr�-  G?��+���uX   DTr�-  j�  �r�-  h h(h
c__builtin__
__main__
hNN}r�-  Ntr�-  Rr�-  �r�-  Rr�-  (X   JJr�-  G?���[�	�X   DTr�-  G?ʐ��[�
X   INr�-  G?���[�	�X   TOr�-  G?�&�9�V�X   VBNr�-  G?���[�	�X   WPr�-  G?�R�+x�X   RBr�-  G?���[�	�X   VBGr�-  G?��+x�5"X   PRPr�-  G?��+x�5"X   PRP$r�-  G?��+x�5"X   RPr�-  G?��+x�5"X   NNr�-  G?�R�+x�X   NNPr�-  G?����[�
hMG?�R�+x�X   NNSr�-  G?��+x�5"X   VBr�-  G?�R�+x�uX   DTr�-  j  �r�-  h h(h
c__builtin__
__main__
hNN}r�-  Ntr�-  Rr�-  �r�-  Rr�-  (X   NNr�-  G?��SIkX   JJr�-  G?�@�z��X   NNSr�-  G?�&�9�V�X   NNPr�-  G?��y��bX   INr�-  G?�@�z�ѡX   CCr�-  G?���<�BX   CDr�-  G?����E�X   VBGr�-  G?�/U�4*�X   VBNr�-  G?�/U�4*�X   WPr�-  G?~���E�hMG?�/U�4*�X   VBDr�-  G?~���E�X   VBr�-  G?~���E�uX   VBPr�-  j�(  �r�-  h h(h
c__builtin__
__main__
hNN}r�-  Ntr�-  Rr�-  �r�-  Rr�-  (X   INr�-  G?�ډ]���X   DTr�-  G?������X   NNPr�-  G?������X   VBNr�-  G?»Q+��X   JJr�-  G?��Q+��X   TOr�-  G?�81�8X   VBGr�-  G?������X   CDr�-  G?������X   RBr�-  G?������X   NNSr�-  G?��Q+��X   RBSr�-  G?������X   PRPr�-  G?������uX   NNPr .  h��r.  h h(h
c__builtin__
__main__
hNN}r.  Ntr.  Rr.  �r.  Rr.  (X   JJr.  G?�E�t]FX   NNr.  G?�]E�t]X   NNSr	.  G?�E�t]FX   NNPr
.  G?�E�t]FuX   INr.  j�  �r.  h h(h
c__builtin__
__main__
hNN}r.  Ntr.  Rr.  �r.  Rr.  (X   NNSr.  G?�������X   NNr.  G?ӻ�����X   INr.  G?�DDDDDDX   NNPr.  G?�333333X   CCr.  G?�UUUUUUh�G?�X   JJr.  G?�UUUUUUX   VBZr.  G?�������X   VBGr.  G?�������X   ``r.  G?�X   VBNr.  G?�X   RBr.  G?�uj�  j.  �r.  h h(h
c__builtin__
__main__
hNN}r.  Ntr.  Rr .  �r!.  Rr".  (X   INr#.  G?��򆼢X   VBDr$.  G?�ה5�yX   MDr%.  G?�ה5�yh�G?̡�(k�X   WPr&.  G?�򆼡�(X   VBNr'.  G?��yC^QX   VBPr(.  G?�(k��X   WRBr).  G?z򆼡�(X   VBZr*.  G?��5�yChMG?�5�yC^X   CCr+.  G?�5�yC^X   VBGr,.  G?�ה5�yX   VBr-.  G?�ה5�yX   TOr..  G?�򆼡�(X   NNSr/.  G?�ה5�yX   JJr0.  G?�򆼡�(NG?�5�yC^X   RBr1.  G?�ה5�yX   WDTr2.  G?z򆼡�(X   ''r3.  G?�5�yC^uX   RBr4.  j   �r5.  h h(h
c__builtin__
__main__
hNN}r6.  Ntr7.  Rr8.  �r9.  Rr:.  (X   VBDr;.  G?��@�´HX   NNr<.  G?�=K��'�h�G?�����]�X   oovr=.  G?��@�´HX   NNPr>.  G?Ţ@�´HX   CCr?.  G?�=K��'�X   POSr@.  G?��V��X   VBNrA.  G?��V��X   WPrB.  G?��V��X   INrC.  G?�9��6X   PRPrD.  G?��V��hMG?��@�´HX   VBrE.  G?�9��6X   VBPrF.  G?��V��X   MDrG.  G?��V��X   NNSrH.  G?��V��X   TOrI.  G?��V��X   RBrJ.  G?��V��X   VBGrK.  G?��V��X   RBSrL.  G?��V��X   JJrM.  G?��@�´HuX   VBDrN.  j�  �rO.  h h(h
c__builtin__
__main__
hNN}rP.  NtrQ.  RrR.  �rS.  RrT.  (X   VBDrU.  G?�      X   NNPrV.  G?�����/hX   NNrW.  G?�q�q�X   RBrX.  G?�����/hX   DTrY.  G?�����/hX   VBrZ.  G?�����/hX   VBNr[.  G?�����/X   VBZr\.  G?�����/hX   JJr].  G?�q�q�X   VBGr^.  G?�q�q�X   WRBr_.  G?�����/hX   oovr`.  G?�����/huj�  j�  �ra.  h h(h
c__builtin__
__main__
hNN}rb.  Ntrc.  Rrd.  �re.  Rrf.  (h�G?��u����X   NNrg.  G?�x��%�X   TOrh.  G?��L�Z��X   INri.  G?��&/5X   VBNrj.  G?�ŀxa�X   NNPrk.  G?�Nl�.�X   WPrl.  G?~s�$}�X   VBGrm.  G?�P�i%njX   DTrn.  G?�_��4J}X   NNSro.  G?��r�`޵X   RPrp.  G?��V�^=X   PRP$rq.  G?��:����X   RBrr.  G?��:����X   WRBrs.  G?��=�X   JJrt.  G?��]K͗X   VBZru.  G?x����X   PRPrv.  G?x����X   VBDrw.  G?b��~�X   VBrx.  G?x����X   oovry.  G?u�L�[X   JJRrz.  G?h����X   CCr{.  G?b��~�X   WDTr|.  G?h����X   MDr}.  G?r��~�X   VBPr~.  G?X����X   NNPSr.  G?b��~�X   ``r�.  G?b��~�hMG?b��~�X   CDr�.  G?X����uX   RBr�.  j�  �r�.  h h(h
c__builtin__
__main__
hNN}r�.  Ntr�.  Rr�.  �r�.  Rr�.  (X   DTr�.  G?�E�t]Fh�G?�E�t]FX   INr�.  G?�t]E�tX   VBZr�.  G?�E�t]Fuj�  j�.  �r�.  h h(h
c__builtin__
__main__
hNN}r�.  Ntr�.  Rr�.  �r�.  Rr�.  (X   NNr�.  G?��LR��&X   NNSr�.  G?���O�X   JJr�.  G?�wA1J��X   NNPr�.  G?���	�VX   VBZr�.  G?yp���rX   JJSr�.  G?�p���rX   CDr�.  G?���	�VX   VBGr�.  G?��6�X   INr�.  G?���	�VX   NNPSr�.  G?�p���rX   DTr�.  G?���	�VX   JJRr�.  G?yp���rX   ``r�.  G?yp���rX   RBSr�.  G?yp���rX   MDr�.  G?yp���rX   oovr�.  G?yp���ruX   TOr�.  j�  �r�.  h h(h
c__builtin__
__main__
hNN}r�.  Ntr�.  Rr�.  �r�.  Rr�.  (h�G?���"��`X   NNPr�.  G?�z�G�{X   NNr�.  G?��O�;dZX   CDr�.  G?�bM���X   NNSr�.  G?�z�G�{hMG?��t�j~�X   DTr�.  G?��t�j~�X   WRBr�.  G?�z�G�{X   VBDr�.  G?��t�j~�X   VBNr�.  G?��t�j~�X   INr�.  G?�bM���X   POSr�.  G?�bM���X   VBr�.  G?�bM���X   JJr�.  G?�bM���NG?�bM���X   WPr�.  G?�z�G�{X   CCr�.  G?�bM���X   VBZr�.  G?�bM���X   oovr�.  G?�bM���uj  j	  �r�.  h h(h
c__builtin__
__main__
hNN}r�.  Ntr�.  Rr�.  �r�.  Rr�.  (X   NNr�.  G?�����X   JJr�.  G?�ƣ�ƣ�X   NNSr�.  G?�恗恘X   NNPr�.  G?æœ�ŔX   VBZr�.  G?y~h~hX   CDr�.  G?�����X   VBNr�.  G?�~h~hX   DTr�.  G?y~h~hX   VBDr�.  G?�^�^�X   NNPSr�.  G?�>�>�X   JJRr�.  G?p����X   INr�.  G?y~h~hX   VBPr�.  G?p����X   VBGr�.  G?�>�>�X   JJSr�.  G?p����X   ``r�.  G?p����uj�+  j�
  �r�.  h h(h
c__builtin__
__main__
hNN}r�.  Ntr�.  Rr�.  �r�.  Rr�.  (X   NNPr�.  G?�q�q�X   INr�.  G?�UUUUUUX   DTr�.  G?�X   VBNr�.  G?��l�lX   WPr�.  G?��l�lX   JJRr�.  G?�X   JJr�.  G?�������X   VBGr�.  G?�X   oovr�.  G?��l�lX   TOr�.  G?�X   NNSr�.  G?�-��-��X   NNr�.  G?�q�q�X   VBr�.  G?��l�lX   RBSr�.  G?�X   PRPr�.  G?��l�lX   RBr�.  G?�������X   PRP$r�.  G?�X   NNPSr�.  G?��l�lX   RPr�.  G?�X   CCr�.  G?�X   ``r�.  G?��l�luX   WDTr�.  j0  �r�.  h h(h
c__builtin__
__main__
hNN}r�.  Ntr�.  Rr�.  �r�.  Rr�.  (X   VBDr�.  G?ڪ�����X   VBZr�.  G?Ҫ�����X   VBPr�.  G?�UUUUUUX   NNSr�.  G?�UUUUUUX   MDr�.  G?�      uj�,  j�&  �r�.  h h(h
c__builtin__
__main__
hNN}r�.  Ntr�.  Rr�.  �r�.  Rr�.  (X   DTr�.  G?�Ye�Ye�X   NNr�.  G?�Ye�Ye�X   NNPr�.  G?�a�a�X   NNSr�.  G?�QEQEX   TOr /  G?�AAX   VBNr/  G?�AAX   CCr/  G?�AAX   INr/  G?�QEQEX   MDr/  G?�AAX   JJr/  G?�a�a�X   ``r/  G?�AAX   WPr/  G?�AAX   PRP$r/  G?�AAX   RPr	/  G?�AAuj�  j\$  �r
/  h h(h
c__builtin__
__main__
hNN}r/  Ntr/  Rr/  �r/  Rr/  (X   RBr/  G?����X   DTr/  G?���*:�X   VBr/  G?ϫ��Tt X   PRPr/  G?����?WX   NNSr/  G?����Tt X   NNPr/  G?�dI囶X   JJr/  G?����X   CDr/  G?����X   NNr/  G?����uj\$  j/  �r/  h h(h
c__builtin__
__main__
hNN}r/  Ntr/  Rr/  �r/  Rr/  (X   VBr/  G?���6�h�G?������X   RBr /  G?������X   NNr!/  G?�ہ�i�X   TOr"/  G?q�|g��X   DTr#/  G?����?X   MDr$/  G?z�:��TX   JJr%/  G?������X   NNPr&/  G?�ہ�i�X   oovr'/  G?��|g��X   VBGr(/  G?q�|g��X   CCr)/  G?q�|g��X   INr*/  G?q�|g��uX   VBNr+/  j  �r,/  h h(h
c__builtin__
__main__
hNN}r-/  Ntr./  Rr//  �r0/  Rr1/  (X   VBDr2/  G?�;�6w�mX   INr3/  G?Ȃ�1rbh�G?Ȃ�1rbX   DTr4/  G?�Ɉ+�WX   MDr5/  G?�W& �LAX   POSr6/  G?�Ɉ+�WX   RBr7/  G?�Ɉ+�WX   ``r8/  G?�Ɉ+�WX   TOr9/  G?�;�6w�mX   JJr:/  G?�Ɉ+�WX   NNr;/  G?�Ɉ+�WX   VBPr</  G?�Ɉ+�WuX   JJr=/  jU  �r>/  h h(h
c__builtin__
__main__
hNN}r?/  Ntr@/  RrA/  �rB/  RrC/  (X   VBDrD/  G?�5�yC^X   NNSrE/  G?�yC^P�X   JJrF/  G?�ה5�yX   VBZrG/  G?��5�yCX   VBPrH/  G?�򆼡�(X   NNPrI/  G?�򆼡�(X   INrJ/  G?��5�yChMG?�򆼡�(X   NNrK/  G?�ה5�yh�G?�5�yC^X   VBGrL/  G?�򆼡�(X   VBNrM/  G?�5�yC^X   CCrN/  G?�5�yC^ujU  jD/  �rO/  h h(h
c__builtin__
__main__
hNN}rP/  NtrQ/  RrR/  �rS/  RrT/  (X   NNPrU/  G?�333333X   DTrV/  G?�333333X   CDrW/  G?ə�����X   TOrX/  G?ə�����uX   NNPrY/  j�  �rZ/  h h(h
c__builtin__
__main__
hNN}r[/  Ntr\/  Rr]/  �r^/  Rr_/  (X   VBDr`/  G?���AI�X   CDra/  G?��.c��X   RBrb/  G?��.c��X   NNrc/  G?�YW��(h�G?�}l=�3�X   VBPrd/  G?����X   VBZre/  G?��:j�pX   JJrf/  G?�}l=�3�X   NNPrg/  G?�}l=�3�X   INrh/  G?�}l=�3�X   MDri/  G?��.c��X   WRBrj/  G?�}l=�3�X   JJRrk/  G?�}l=�3�X   NNSrl/  G?�}l=�3�uX   PRPrm/  j�  �rn/  h h(h
c__builtin__
__main__
hNN}ro/  Ntrp/  Rrq/  �rr/  Rrs/  (h�G?��;�6xX   DTrt/  G?�;�6w�mX   INru/  G?�W& �LX   TOrv/  G?�W& �LX   NNPrw/  G?�Ɉ+�WX   WDTrx/  G?�Ɉ+�WX   NNry/  G?�W& �LAX   JJrz/  G?�Ɉ+�WX   VBNr{/  G?�W& �LAX   RBr|/  G?�W& �LAX   WRBr}/  G?�Ɉ+�Wuj�+  j  �r~/  h h(h
c__builtin__
__main__
hNN}r/  Ntr�/  Rr�/  �r�/  Rr�/  (h�G?�|�`�g�X   NNSr�/  G?�7Y�)�vX   INr�/  G?���ϑLhMG?���ϑLX   WPr�/  G?������X   VBDr�/  G?���ϑLX   WRBr�/  G?������X   NNr�/  G?���ϑLX   VBNr�/  G?������X   VBGr�/  G?������X   RBr�/  G?������X   ''r�/  G?������X   POSr�/  G?������X   TOr�/  G?������uX   PRP$r�/  j�  �r�/  h h(h
c__builtin__
__main__
hNN}r�/  Ntr�/  Rr�/  �r�/  Rr�/  (X   NNr�/  G?ډ]��ډX   JJr�/  G?��Q+��X   VBNr�/  G?������X   DTr�/  G?������X   WPr�/  G?������X   RBr�/  G?������X   NNSr�/  G?�ډ]���X   INr�/  G?������X   NNPr�/  G?������uX   VBPr�/  j�  �r�/  h h(h
c__builtin__
__main__
hNN}r�/  Ntr�/  Rr�/  �r�/  Rr�/  (X   NNSr�/  G?�WWWWWWX   INr�/  G?ٙ�����X   JJr�/  G?�X   VBr�/  G?�X   NNr�/  G?�h�G?�X   CDr�/  G?�X   TOr�/  G?�X   CCr�/  G?�uX   oovr�/  j�  �r�/  h h(h
c__builtin__
__main__
hNN}r�/  Ntr�/  Rr�/  �r�/  Rr�/  (X   VBDr�/  G?�I���T�X   INr�/  G?Ϫ�I��h�G?�;���X   NNr�/  G?�����X   oovr�/  G?����X   TOr�/  G?����X   NNSr�/  G?�{y�!��X   CCr�/  G?������X   WRBr�/  G?�I���T�X   WPr�/  G?q���X   VBGr�/  G?�I���T�X   VBPr�/  G?����hMG?������X   JJr�/  G?�(�5�2�NG?q���X   NNPr�/  G?������X   VBNr�/  G?y�����X   VBZr�/  G?q���X   RBr�/  G?y�����X   DTr�/  G?q���X   ``r�/  G?q���uX   POSr�/  h��r�/  h h(h
c__builtin__
__main__
hNN}r�/  Ntr�/  Rr�/  �r�/  Rr�/  NG?�      sX   VBDr�/  j�  �r�/  h h(h
c__builtin__
__main__
hNN}r�/  Ntr�/  Rr�/  �r�/  Rr�/  (h�G?�&ɲl�'X   NNSr�/  G?�d�6M�eX   NNr�/  G?�      X   NNPr�/  G?���|X   INr�/  G?�l�&ɲmX   JJr�/  G?�6M�d�6X   TOr�/  G?�&ɲl�'X   VBNr�/  G?�E�t]FX   VBGr�/  G?�E�t]FX   RBr�/  G?���|X   VBr�/  G?���|uj�  h��r�/  h h(h
c__builtin__
__main__
hNN}r�/  Ntr�/  Rr�/  �r�/  Rr�/  NG?�      sX   JJr�/  j  �r�/  h h(h
c__builtin__
__main__
hNN}r�/  Ntr�/  Rr�/  �r�/  Rr�/  (X   VBDr�/  G?�A�A�X   MDr�/  G?��_�_X   VBZr�/  G?ə�����hMG?�A�A�X   VBPr�/  G?�A�A�X   NNSr�/  G?�A�A�X   JJr�/  G?�A�A�X   INr�/  G?ə�����X   oovr�/  G?�A�A�X   ``r�/  G?�A�A�uX   CCr�/  j�  �r�/  h h(h
c__builtin__
__main__
hNN}r�/  Ntr�/  Rr�/  �r�/  Rr�/  (X   NNSr�/  G?�)�B�X   NNr�/  G?һQ+��h�G?����X   RBr�/  G?���
h�X   WPr 0  G?���
h�X   INr0  G?������X   VBGr0  G?���
h�X   WRBr0  G?���
h�X   JJr0  G?������X   VBNr0  G?���
h�X   JJRr0  G?���
h�X   VBDr0  G?���
h�X   TOr0  G?������hMG?���
h�uX   NNPr	0  h��r
0  h h(h
c__builtin__
__main__
hNN}r0  Ntr0  Rr0  �r0  Rr0  (X   oovr0  G?��h`��CX   NNPr0  G?ןP4���X   CDr0  G?�����l�X   RBr0  G?����>X   DTr0  G?��L��RgX   CCr0  G?����6�h�G?�S����X   JJr0  G?��S����X   VBPr0  G?�^}@���X   NNr0  G?�����mX   VBDr0  G?����6�X   NNSr0  G?��#(�X   INr0  G?�+���_�X   VBZr0  G?��S����X   VBr0  G?�Ò ��X   PRPr0  G?q�S����X   VBNr0  G?��S����hMG?q�S����X   ''r 0  G?q�S����NG?q�S����X   NNPSr!0  G?q�S����X   WPr"0  G?z^}@���X   JJSr#0  G?q�S����X   VBGr$0  G?q�S����X   WRBr%0  G?z^}@���X   ``r&0  G?q�S����uh�j0  �r'0  h h(h
c__builtin__
__main__
hNN}r(0  Ntr)0  Rr*0  �r+0  Rr,0  (X   oovr-0  G?Ƶ�kZֶX   VBNr.0  G?��!B�h�G?��!B�X   JJr/0  G?��!B�X   NNPr00  G?Є!B�X   NNr10  G?Ƶ�kZֶX   TOr20  G?��1�c�X   VBGr30  G?��!B�X   DTr40  G?��!B�X   VBPr50  G?��!B�X   CDr60  G?��1�c�X   ``r70  G?��!B�uX   NNSr80  j[)  �r90  h h(h
c__builtin__
__main__
hNN}r:0  Ntr;0  Rr<0  �r=0  Rr>0  (X   INr?0  G?��9Z��ph�G?��<'+]�X   RBr@0  G?�ƥ/�X   TOrA0  G?��g��k�X   VBDrB0  G?��0�5)X   VBPrC0  G?�|��cSX   CCrD0  G?�/�a�jX   VBNrE0  G?��ͣ��X   MDrF0  G?��qO��;X   WPrG0  G?��g��k�X   WDTrH0  G?��qO��;X   VBGrI0  G?������X   NNrJ0  G?��qO��;X   DTrK0  G?va�jQ"�X   CDrL0  G?va�jQ"�X   VBZrM0  G?��g��k�hMG?��g��k�X   NNPrN0  G?��g��k�NG?va�jQ"�X   VBrO0  G?�a�jQ"�X   NNSrP0  G?�a�jQ"�X   RBSrQ0  G?va�jQ"�X   JJrR0  G?��qO��;X   WRBrS0  G?va�jQ"�X   JJRrT0  G?va�jQ"�uX   oovrU0  h��rV0  h h(h
c__builtin__
__main__
hNN}rW0  NtrX0  RrY0  �rZ0  Rr[0  (NG?��<��<�h�G?�y�y�X   ''r\0  G?�I$�I$�hMG?�I$�I$�uX   VBNr]0  j+!  �r^0  h h(h
c__builtin__
__main__
hNN}r_0  Ntr`0  Rra0  �rb0  Rrc0  (X   NNPrd0  G?س�,�:X   JJre0  G?�ה5�yX   NNrf0  G?�򆼡�(X   INrg0  G?��}�pX   DTrh0  G?�򆼡�(X   JJRri0  G?�򆼡�(h�G?�򆼡�(uX   ''rj0  j�  �rk0  h h(h
c__builtin__
__main__
hNN}rl0  Ntrm0  Rrn0  �ro0  Rrp0  (h�G?ٰ�6X   INrq0  G?ٰ�6X   TOrr0  G?�Ի~2z�X   RBrs0  G?��@�´HX   NNSrt0  G?��@�´HX   VBNru0  G?��V��X   DTrv0  G?��V��X   RPrw0  G?��V��X   ``rx0  G?��@�´HuX   VBry0  j,  �rz0  h h(h
c__builtin__
__main__
hNN}r{0  Ntr|0  Rr}0  �r~0  Rr0  (X   NNPr�0  G?���n�X   VBr�0  G?��1�c�X   NNSr�0  G?��!B�X   RBr�0  G?��`XX   NNr�0  G?���n�X   TOr�0  G?��`XX   VBGr�0  G?��!B�X   JJr�0  G?���n�X   VBDr�0  G?��!B�X   VBPr�0  G?��`XX   INr�0  G?��`XX   WPr�0  G?��!B�X   MDr�0  G?��`XuX   NNSr�0  j�  �r�0  h h(h
c__builtin__
__main__
hNN}r�0  Ntr�0  Rr�0  �r�0  Rr�0  (X   NNr�0  G?�&	��hX   JJr�0  G?�"���b*X   NNSr�0  G?�R�T�,X   VBPr�0  G?�����X   JJSr�0  G?~����X   VBZr�0  G?~����X   INr�0  G?�����X   NNPr�0  G?��Aq�X   VBGr�0  G?��Aq�X   ``r�0  G?�?���3�X   VBNr�0  G?�?���3�X   TOr�0  G?��Aq�h�G?�,EKR�X   VBDr�0  G?~����X   DTr�0  G?~����X   CCr�0  G?~����X   RBr�0  G?��Aq�uNh-�r�0  h h(h
c__builtin__
__main__
hNN}r�0  Ntr�0  Rr�0  �r�0  Rr�0  (X   VBPr�0  G?��t]E�X   DTr�0  G?�t]E�tX   VBZr�0  G?��t]E�X   INr�0  G?�E�t]FX   NNSr�0  G?�E�t]FX   NNPr�0  G?�E�t]FX   CDr�0  G?�]E�t]X   RBr�0  G?�E�t]FX   VBDr�0  G?�E�t]FX   JJr�0  G?�E�t]FX   MDr�0  G?�E�t]FX   WPr�0  G?�E�t]Fuh-j�0  �r�0  h h(h
c__builtin__
__main__
hNN}r�0  Ntr�0  Rr�0  �r�0  Rr�0  (X   INr�0  G?���J3�)X   CDr�0  G?�B�Y!dX   JJr�0  G?��`v���X   VBNr�0  G?���J3�)X   RBr�0  G?�B�Y!dX   DTr�0  G?��`v��X   NNSr�0  G?�B�Y!dX   JJRr�0  G?���J3�)X   VBZr�0  G?��`v���X   RPr�0  G?��`v���X   WRBr�0  G?�B�Y!dX   TOr�0  G?�B�Y!dX   VBGr�0  G?��`v���h�G?�B�Y!duX   VBGr�0  j}  �r�0  h h(h
c__builtin__
__main__
hNN}r�0  Ntr�0  Rr�0  �r�0  Rr�0  (X   NNr�0  G?ܰ�=��X   VBZr�0  G?�{���aX   NNPr�0  G?�{���aX   CDr�0  G?���a{�X   NNSr�0  G?�{���aX   JJr�0  G?�{���aX   VBDr�0  G?���a{�uj	  j
!  �r�0  h h(h
c__builtin__
__main__
hNN}r�0  Ntr�0  Rr�0  �r�0  Rr�0  (X   VBr�0  G?��t�j~�h�G?θQ��X   DTr�0  G?�bM���X   VBZr�0  G?�z�G�{X   JJr�0  G?�bM���X   TOr�0  G?��+I�X   VBPr�0  G?�bM���X   INr�0  G?Ͼvȴ9XhMG?�bM���X   MDr�0  G?��t�j~�X   RBr�0  G?�bM���X   WPr�0  G?�bM���X   ''r�0  G?�bM���X   CDr�0  G?�bM���X   VBDr�0  G?��t�j~�X   PRP$r�0  G?�bM���X   CCr�0  G?�bM���X   RPr�0  G?�bM���X   NNr�0  G?��t�j~�X   WRBr�0  G?�bM���X   ``r�0  G?��t�j~�uj�0  hM�r�0  h h(h
c__builtin__
__main__
hNN}r�0  Ntr�0  Rr�0  �r�0  Rr�0  (X   WPr�0  G?�yf톙X   JJr�0  G?����Tt X   VBGr�0  G?�yf톙X   WDTr�0  G?����X   NNPr�0  G?����X   INr�0  G?�dI囶X   oovr�0  G?����Tt X   ''r�0  G?����X   VBr�0  G?����X   NNr�0  G?����Tt X   DTr 1  G?�dI囶X   CCr1  G?����Tt X   RBr1  G?����X   PRPr1  G?����X   VBNr1  G?����Tt X   JJSr1  G?����X   VBZr1  G?����X   NNSr1  G?����Tt X   WRBr1  G?����X   ``r	1  G?����uj�  j�  �r
1  h h(h
c__builtin__
__main__
hNN}r1  Ntr1  Rr1  �r1  Rr1  (X   MDr1  G?�������X   JJr1  G?�333333X   NNr1  G?�      X   NNSr1  G?ə�����X   NNPr1  G?�������uj�  j1  �r1  h h(h
c__builtin__
__main__
hNN}r1  Ntr1  Rr1  �r1  Rr1  (h�G?�      X   INr1  G?�      X   VBNr1  G?�      X   CCr1  G?�      uj1  h��r1  h h(h
c__builtin__
__main__
hNN}r1  Ntr 1  Rr!1  �r"1  Rr#1  NG?�      sj�  hc�r$1  h h(h
c__builtin__
__main__
hNN}r%1  Ntr&1  Rr'1  �r(1  Rr)1  (X   PRPr*1  G?�A�A�X   CDr+1  G?��;�;X   RBr,1  G?��;�;X   DTr-1  G?�i�i�X   INr.1  G?�i�i�X   VBr/1  G?�A�A�X   JJr01  G?��;�;X   NNSr11  G?�A�A�X   NNPr21  G?�A�A�X   NNr31  G?��;�;uhMj0  �r41  h h(h
c__builtin__
__main__
hNN}r51  Ntr61  Rr71  �r81  Rr91  (X   JJr:1  G?��;�;X   NNr;1  G?��y���hMG?̤�^�X   MDr<1  G?|��^�X   VBNr=1  G?���^�X   INr>1  G?��;�;X   NNSr?1  G?��>�G��X   CCr@1  G?��K0U�X   NNPrA1  G?����[L�h�G?���^�X   VBGrB1  G?|��^�X   TOrC1  G?�{�D)-X   CDrD1  G?|��^�uX   VBPrE1  j�  �rF1  h h(h
c__builtin__
__main__
hNN}rG1  NtrH1  RrI1  �rJ1  RrK1  (X   INrL1  G?�$l+D�X   JJrM1  G?�=K��'�X   RPrN1  G?��V��X   NNSrO1  G?ό����X   NNrP1  G?Ļ~2z�pX   VBrQ1  G?��V��X   CCrR1  G?��@�´HX   TOrS1  G?�6�@�X   VBGrT1  G?��V��X   VBNrU1  G?��V��X   NNPrV1  G?��V��hMG?��V��X   RBrW1  G?��V��X   VBZrX1  G?��V��X   WPrY1  G?��V��uj�  jL1  �rZ1  h h(h
c__builtin__
__main__
hNN}r[1  Ntr\1  Rr]1  �r^1  Rr_1  (X   DTr`1  G?̏#��<�X   NNSra1  G?�e�v]�fX   WPrb1  G?��yG��X   VBGrc1  G?��1�c�X   CDrd1  G?�����{�X   WRBre1  G?��!B�X   NNPrf1  G?�G��yHX   VBNrg1  G?���n�X   NNrh1  G?�UUUUUUX   INri1  G?��!B�X   oovrj1  G?��!B�X   JJrk1  G?�D�4MEX   RBrl1  G?���n�X   PRPrm1  G?��1�c�h�G?��!B�X   PRP$rn1  G?��1�c�X   JJSro1  G?���n�X   TOrp1  G?��!B�X   WDTrq1  G?v�`XX   JJRrr1  G?��!B�X   ``rs1  G?v�`XX   CCrt1  G?v�`Xuj�"  j�'  �ru1  h h(h
c__builtin__
__main__
hNN}rv1  Ntrw1  Rrx1  �ry1  Rrz1  (X   WPr{1  G?��\��X   VBNr|1  G?�o��,bGX   NNSr}1  G?���	��X   RBr~1  G?�f=���X   JJr1  G?��d�W/X   VBr�1  G?��Rm_�X   VBDr�1  G?��r!I��X   DTr�1  G?��r!I��X   NNPr�1  G?���}9�X   PRP$r�1  G?��ڿ�F�X   NNr�1  G? \��X   VBGr�1  G?�����U�X   JJRr�1  G?����U�X   NNPSr�1  G?y\��w�X   VBZr�1  G?�򆼡�(X   WDTr�1  G?i\��w�X   INr�1  G?|�Rm_�X   CDr�1  G?����U�X   TOr�1  G?Y\��w�X   VBPr�1  G?|�Rm_�X   JJSr�1  G?o����U�X   WRBr�1  G?y\��w�X   oovr�1  G?c�H��X   ``r�1  G?Y\��w�X   PRPr�1  G?c�H��X   MDr�1  G?Y\��w�X   CCr�1  G?Y\��w�uX   CDr�1  j_  �r�1  h h(h
c__builtin__
__main__
hNN}r�1  Ntr�1  Rr�1  �r�1  Rr�1  (X   JJr�1  G?�<<<<<<X   NNSr�1  G?�uX   WPr�1  jZ%  �r�1  h h(h
c__builtin__
__main__
hNN}r�1  Ntr�1  Rr�1  �r�1  Rr�1  (X   RBr�1  G?�      X   INr�1  G?�      X   VBPr�1  G?�      X   VBZr�1  G?�      X   VBDr�1  G?�      X   JJr�1  G?�      ujZ%  j�1  �r�1  h h(h
c__builtin__
__main__
hNN}r�1  Ntr�1  Rr�1  �r�1  Rr�1  (X   VBNr�1  G?����:�X   RBr�1  G?�ȿ�!'X   JJr�1  G?�w�T�,4X   INr�1  G?�V����X   oovr�1  G?�w�T�,4h�G?�ȿ�!&�X   VBr�1  G?��V����X   VBDr�1  G?�w�T�,4X   DTr�1  G?�j����X   JJRr�1  G?�ȿ�!'X   VBZr�1  G?�ȿ�!'X   TOr�1  G?�w�T�,4X   VBPr�1  G?�w�T�,4X   CCr�1  G?�w�T�,4X   NNPr�1  G?�ȿ�!'hMG?�w�T�,4X   NNSr�1  G?�w�T�,4X   VBGr�1  G?�ȿ�!'uX   VBNr�1  j  �r�1  h h(h
c__builtin__
__main__
hNN}r�1  Ntr�1  Rr�1  �r�1  Rr�1  (X   INr�1  G?�W& �LX   NNr�1  G?�W& �Lh�G?�Ɉ+�WX   NNSr�1  G?�W& �LAX   JJr�1  G?�W& �LAX   TOr�1  G?�W& �LAX   RBr�1  G?�Ɉ+�WX   CCr�1  G?�Ɉ+�WX   WPr�1  G?�Ɉ+�WuX   CDr�1  j�
  �r�1  h h(h
c__builtin__
__main__
hNN}r�1  Ntr�1  Rr�1  �r�1  Rr�1  (X   NNr�1  G?�a�a�X   NNSr�1  G?�a�a�X   INr�1  G?�I$�I$�X   PRP$r�1  G?�a�a�X   JJr�1  G?�a�a�h�G?�a�a�X   NNPr�1  G?�a�a�uX   VBPr�1  jL  �r�1  h h(h
c__builtin__
__main__
hNN}r�1  Ntr�1  Rr�1  �r�1  Rr�1  (X   VBNr�1  G?�0�_��X   TOr�1  G?�	���`X   INr�1  G?�K�3��HX   VBr�1  G?��{.oNX   RBr�1  G?��Ҟ�jX   VBGr�1  G?�;f�PmWX   VBPr�1  G?�9]d��X   JJr�1  G?�Sg�+t�X   WPr�1  G?��DV5�:h�G?�X�x�K,X   WDTr�1  G?��A���X   CCr�1  G?���d��CX   VBDr�1  G?��Ҟ�jhMG?|	���`X   VBZr�1  G?l	���`X   NNSr�1  G?��DV5�:X   POSr�1  G?�	���`X   MDr�1  G?`�DV5�:X   NNPr�1  G?s��d��CX   WRBr�1  G?Vm�r�(MX   oovr�1  G?Vm�r�(MX   DTr�1  G?`�DV5�:X   RBSr�1  G?fm�r�(MX   NNr�1  G?s��d��CNG?Vm�r�(MX   JJRr�1  G?`�DV5�:X   ''r�1  G?Vm�r�(MX   CDr�1  G?Vm�r�(MX   ``r�1  G?Vm�r�(MuX   INr�1  jI  �r 2  h h(h
c__builtin__
__main__
hNN}r2  Ntr2  Rr2  �r2  Rr2  (X   NNSr2  G?������X   DTr2  G?������h�G?�����hMG?������X   PRP$r2  G?������X   PRPr	2  G?��Q+��X   TOr
2  G?������X   JJr2  G?��Q+��X   WRBr2  G?������X   NNr2  G?������X   RPr2  G?������X   NNPr2  G?������uX   NNr2  j   �r2  h h(h
c__builtin__
__main__
hNN}r2  Ntr2  Rr2  �r2  Rr2  (X   INr2  G?�h�G?�ZZZZZZX   VBr2  G?�X   CCr2  G?�������X   NNr2  G?�ZZZZZZX   RPr2  G?�X   NNSr2  G?�������X   VBDr2  G?�X   MDr2  G?�X   JJr2  G?�uX   CCr 2  j�  �r!2  h h(h
c__builtin__
__main__
hNN}r"2  Ntr#2  Rr$2  �r%2  Rr&2  (X   INr'2  G?�cp!���X   DTr(2  G?�
�cp"X   TOr)2  G?�cp!���X   PRP$r*2  G?���k朐X   JJr+2  G?�cp!���X   VBNr,2  G?���V�jX   RBr-2  G?���|ӑ�X   NNPr.2  G?�(2��C�X   NNr/2  G?���k朐X   RPr02  G?�(2��C�X   PRPr12  G?���|ӑ�X   NNSr22  G?���k朐X   JJRr32  G?���k朐X   oovr42  G?���k朐X   RBSr52  G?���k朐X   JJSr62  G?�cp!���X   VBGr72  G?���k朐X   CDr82  G?���k朐uX   VBZr92  jN  �r:2  h h(h
c__builtin__
__main__
hNN}r;2  Ntr<2  Rr=2  �r>2  Rr?2  (X   JJr@2  G?�������X   NNrA2  G?��8�9X   VBDrB2  G?�q�q�X   VBrC2  G?��8�9X   NNSrD2  G?��8�9X   INrE2  G?�8�8�X   NNPrF2  G?��q�rX   RBrG2  G?�UUUUUUhMG?��8�9X   TOrH2  G?�q�q�X   CCrI2  G?�q�q�h�G?��8�9X   CDrJ2  G?�q�q�X   DTrK2  G?�q�q�X   oovrL2  G?�q�q�uX   CDrM2  jl-  �rN2  h h(h
c__builtin__
__main__
hNN}rO2  NtrP2  RrQ2  �rR2  RrS2  (X   DTrT2  G?�A�A�X   INrU2  G?ə�����X   VBNrV2  G?�A�A�X   RBrW2  G?�I$�I$�X   JJrX2  G?��_�_X   NNSrY2  G?�A�A�h�G?�A�A�NG?�A�A�X   PRPrZ2  G?�A�A�X   oovr[2  G?�A�A�ujJ  j  �r\2  h h(h
c__builtin__
__main__
hNN}r]2  Ntr^2  Rr_2  �r`2  Rra2  (X   INrb2  G?��_�pr�X   NNrc2  G?Ո_�pr�X   JJrd2  G?��f�宧X   NNSre2  G?�&GƔV!X   ''rf2  G?�#�J+�h�G?�#�J+�X   WPrg2  G?����@�X   CCrh2  G?�#�J+�X   CDri2  G?������X   NNPrj2  G?������hMG?����@�uX   NNSrk2  j�  �rl2  h h(h
c__builtin__
__main__
hNN}rm2  Ntrn2  Rro2  �rp2  Rrq2  (X   TOrr2  G?���7]8OX   INrs2  G?��D��X   NNrt2  G?�E�akjX   VBDru2  G?��nAM"h�G?����	�X   NNSrv2  G?����	�hMG?���N�X   JJrw2  G?����f�X   VBPrx2  G?��nAM"X   VBZry2  G?��nAM"X   CCrz2  G?��5x�Y�X   NNPr{2  G?���N�X   RBr|2  G?����f�X   WRBr}2  G?�틗�=X   VBNr~2  G?v���f�X   DTr2  G?v���f�X   NNPSr�2  G?~H�Yo3�X   VBr�2  G?~H�Yo3�X   VBGr�2  G?nH�Yo3�NG?nH�Yo3�X   JJSr�2  G?nH�Yo3�X   oovr�2  G?nH�Yo3�uj�  j�  �r�2  h h(h
c__builtin__
__main__
hNN}r�2  Ntr�2  Rr�2  �r�2  Rr�2  (X   NNPr�2  G?�UUUUUUX   JJr�2  G?�UUUUUUX   NNr�2  G?�UUUUUUuX   POSr�2  jX  �r�2  h h(h
c__builtin__
__main__
hNN}r�2  Ntr�2  Rr�2  �r�2  Rr�2  (X   NNPr�2  G?�z�G�{X   VBNr�2  G?�
=p��
X   RBr�2  G?�z�G�{X   JJr�2  G?�z�G�{X   DTr�2  G?�������X   VBGr�2  G?�z�G�{X   INr�2  G?�z�G�{X   NNSr�2  G?�z�G�{X   NNPSr�2  G?�z�G�{X   PRPr�2  G?�z�G�{h�G?�z�G�{X   TOr�2  G?�z�G�{uX   NNSr�2  j�  �r�2  h h(h
c__builtin__
__main__
hNN}r�2  Ntr�2  Rr�2  �r�2  Rr�2  (X   INr�2  G?��f�fh�G?�B�B�X   NNr�2  G?��k�kX   VBDr�2  G?�l�l�X   VBNr�2  G?�l�l�X   VBPr�2  G?�g�g�X   DTr�2  G?��p�pX   VBZr�2  G?��p�pX   CCr�2  G?�X   VBr�2  G?��p�pX   RBr�2  G?�X   VBGr�2  G?��p�pX   NNSr�2  G?��f�fX   TOr�2  G?��p�pX   WDTr�2  G?�NG?��p�puX   POSr�2  jY  �r�2  h h(h
c__builtin__
__main__
hNN}r�2  Ntr�2  Rr�2  �r�2  Rr�2  (h�G?��q�rX   VBZr�2  G?�q�q�X   NNPr�2  G?�q�q�uX   WRBr�2  j�  �r�2  h h(h
c__builtin__
__main__
hNN}r�2  Ntr�2  Rr�2  �r�2  Rr�2  (X   INr�2  G?�?]�<��h�G?�F�eb��X   NNSr�2  G?�jt�F�X   TOr�2  G?�F�eb�X   RBr�2  G?�F�eb��X   NNr�2  G?�X�~��zhMG?�jt�F�X   JJr�2  G?�F�eb��X   DTr�2  G?�F�eb��X   RPr�2  G?�F�eb��X   VBZr�2  G?�F�eb��uX   PRPr�2  hM�r�2  h h(h
c__builtin__
__main__
hNN}r�2  Ntr�2  Rr�2  �r�2  Rr�2  (X   VBDr�2  G?�������X   WPr�2  G?�X   INr�2  G?Ɩ�����X   WRBr�2  G?�������X   NNPr�2  G?�X   CCr�2  G?�������X   VBGr�2  G?�h�G?�X   ``r�2  G?�������uX   VBPr�2  j�  �r�2  h h(h
c__builtin__
__main__
hNN}r�2  Ntr�2  Rr�2  �r�2  Rr�2  (X   VBNr�2  G?�[O[OX   JJr�2  G?��$�$X   VBr�2  G?��$�$h�G?�/�/�X   RBr�2  G?�)Z)ZX   INr�2  G?�G�G�X   TOr�2  G?�X   DTr�2  G?�����X   VBGr�2  G?�PPX   WRBr�2  G?^����X   WPr�2  G?��`�`X   NNPr�2  G?�PPX   JJRr�2  G?v�`�`X   NNSr�2  G?�����X   oovr�2  G?�����X   CDr�2  G?�5�5�X   VBDr�2  G?f�`�`X   NNr�2  G?�5�5�X   CCr�2  G?sPPNG?^����X   PRPr�2  G?n����hMG?^����X   VBZr�2  G?^����X   PRP$r�2  G?^����uX   JJr�2  j�   �r�2  h h(h
c__builtin__
__main__
hNN}r�2  Ntr�2  Rr�2  �r�2  Rr�2  (X   NNSr 3  G?�m��m��X   JJSr3  G?�I$�I$�X   NNr3  G?�I$�I$�uX   DTr3  j�  �r3  h h(h
c__builtin__
__main__
hNN}r3  Ntr3  Rr3  �r3  Rr	3  (X   VBDr
3  G?�ʸ�%�X   NNr3  G?���WX   CCr3  G?���Ξ�X   VBGr3  G?�0ʸ�&X   VBr3  G?����X   NNPSr3  G?�1av@��h�G?ɪ;�҄�X   INr3  G?�g����mX   MDr3  G?������8X   NNPr3  G?�J1avAX   VBPr3  G?ç�o���X   WDTr3  G?y�f��JX   PRPr3  G?dʸ�%�nX   ''r3  G?o0ʸ�&X   NNSr3  G?�ʸ�%�nX   JJr3  G?�d�
eX   RBr3  G?��f��JX   WPr3  G?�d�
e\X   TOr3  G?�ʸ�%�nhMG?������8X   VBNr3  G?�1av@��X   DTr3  G?�1av@��X   ``r3  G?0ʸ�&X   WRBr3  G?dʸ�%�nX   VBZr 3  G?0ʸ�&NG?o0ʸ�&X   POSr!3  G?0ʸ�&uj�  j
3  �r"3  h h(h
c__builtin__
__main__
hNN}r#3  Ntr$3  Rr%3  �r&3  Rr'3  (X   INr(3  G?��H���X   VBNr)3  G?�,bGT�h�G?��	��$uX   NNPr*3  G?�򆼡�(X   DTr+3  G?��Rm_�X   RBr,3  G?�X   CDr-3  G?�\��w�X   NNr.3  G?�\��w�X   TOr/3  G?�����U�X   JJSr03  G?�����U�X   JJr13  G?�\��w�X   RBSr23  G?y\��w�X   PRP$r33  G?�����U�X   VBDr43  G?��H��X   VBGr53  G?�\��w�X   VBr63  G?��H��X   WRBr73  G?��H��X   WPr83  G?��Rm_�X   RPr93  G?��H��X   NNSr:3  G?��H��X   WDTr;3  G?��H��NG?��H��X   ``r<3  G?y\��w�X   PRPr=3  G?��H��uX   oovr>3  j�  �r?3  h h(h
c__builtin__
__main__
hNN}r@3  NtrA3  RrB3  �rC3  RrD3  (X   JJrE3  G?��V��X   NNSrF3  G?��V��X   VBrG3  G?�6�@�X   CCrH3  G?��@�´HX   PRPrI3  G?�9��6X   NNPrJ3  G?�=K��'�X   INrK3  G?�6�@�X   DTrL3  G?�6�@�h�G?��V��X   TOrM3  G?��V��X   oovrN3  G?��V��X   RBrO3  G?��@�´HX   VBPrP3  G?��V��X   CDrQ3  G?��V��X   WPrR3  G?��V��X   PRP$rS3  G?��V��X   NNrT3  G?��@�´HX   WRBrU3  G?��V��uj�+  j�  �rV3  h h(h
c__builtin__
__main__
hNN}rW3  NtrX3  RrY3  �rZ3  Rr[3  (X   VBDr\3  G?���a|X   VBZr]3  G?�{���aX   MDr^3  G?�{���aX   VBPr_3  G?�ܰ�=�	X   JJr`3  G?���a{�X   VBra3  G?�{���aX   INrb3  G?���a{�X   NNSrc3  G?���a{�uX   NNPrd3  j�  �re3  h h(h
c__builtin__
__main__
hNN}rf3  Ntrg3  Rrh3  �ri3  Rrj3  (X   NNrk3  G?�������X   DTrl3  G?�X   VBDrm3  G?�h�G?�X   NNSrn3  G?�X   JJro3  G?�X   NNPrp3  G?�X   TOrq3  G?�X   VBNrr3  G?Ɩ�����X   INrs3  G?�X   RBrt3  G?�X   VBru3  G?�NG?�uX   NNPSrv3  j  �rw3  h h(h
c__builtin__
__main__
hNN}rx3  Ntry3  Rrz3  �r{3  Rr|3  (X   NNPr}3  G?ѧ�a{�X   WPr~3  G?��L�x��X   NNPSr3  G?��f��pX   NNSr�3  G?��L�x��X   DTr�3  G?ǊL�x��X   VBDr�3  G?���a{�X   JJr�3  G?���I�/X   PRP$r�3  G?��L�x��uX   VBPr�3  j
  �r�3  h h(h
c__builtin__
__main__
hNN}r�3  Ntr�3  Rr�3  �r�3  Rr�3  (X   TOr�3  G?�{���aX   DTr�3  G?��,#Or�X   VBNr�3  G?���a|X   VBGr�3  G?���a{�X   NNSr�3  G?�{���aX   JJr�3  G?���a{�X   RBr�3  G?�ܰ�=�	X   oovr�3  G?�{���aX   INr�3  G?���a{�X   NNPr�3  G?���a|X   WDTr�3  G?���a{�X   WRBr�3  G?���a{�X   NNr�3  G?�{���aX   RBSr�3  G?���a{�X   PRPr�3  G?���a{�X   JJRr�3  G?�{���ah�G?���a{�X   RPr�3  G?���a{�X   ``r�3  G?�{���auX   NNPSr�3  j  �r�3  h h(h
c__builtin__
__main__
hNN}r�3  Ntr�3  Rr�3  �r�3  Rr�3  (h�G?�W�x�XX   NNPr�3  G?��Y/��X   CCr�3  G?�m��mX   NNr�3  G?�m��mX   VBDr�3  G?���=�X   POSr�3  G?�m��mX   VBNr�3  G?��!B�X   INr�3  G?��!B�X   TOr�3  G?���=�X   VBZr�3  G?�m��mX   WPr�3  G?���=�hMG?���=�X   VBPr�3  G?�m��mX   NNSr�3  G?�m��mX   VBGr�3  G?���=�X   CDr�3  G?���=�X   VBr�3  G?�m��mX   RBr�3  G?�m��mX   NNPSr�3  G?���=�X   ``r�3  G?�m��muj�  j1  �r�3  h h(h
c__builtin__
__main__
hNN}r�3  Ntr�3  Rr�3  �r�3  Rr�3  (X   PRPr�3  G?�UUUUUUX   NNPr�3  G?ʪ�����X   WPr�3  G?�UUUUUUX   NNr�3  G?�UUUUUUX   DTr�3  G?�UUUUUUX   VBNr�3  G?�UUUUUUX   JJSr�3  G?�UUUUUUX   JJr�3  G?�      uX   JJr�3  j�  �r�3  h h(h
c__builtin__
__main__
hNN}r�3  Ntr�3  Rr�3  �r�3  Rr�3  (X   INr�3  G?����� X   DTr�3  G?ڕ�Z��[X   VBr�3  G?ӱ;�;X   JJr�3  G?��z�zX   NNPr�3  G?����� X   PRPr�3  G?��z�zX   NNSr�3  G?����� X   ``r�3  G?����� X   CCr�3  G?����� uj�
  j+  �r�3  h h(h
c__builtin__
__main__
hNN}r�3  Ntr�3  Rr�3  �r�3  Rr�3  (X   VBDr�3  G?���/9X   NNr�3  G?����/NG?���/9X   INr�3  G?�X��ƈX   VBNr�3  G?�I$�I$�X   DTr�3  G?×����X   PRP$r�3  G?���/9h�G?×����X   TOr�3  G?�X��Ƈ�X   NNSr�3  G?�X��Ƈ�X   JJr�3  G?�X��Ƈ�X   VBGr�3  G?���/9X   WPr�3  G?���/9X   NNPr�3  G?���/9uj�  jC  �r�3  h h(h
c__builtin__
__main__
hNN}r�3  Ntr�3  Rr�3  �r�3  Rr�3  (X   NNr�3  G?��zoM�X   JJr�3  G?�B�Y!dX   NNPr�3  G?��zoM�X   VBNr�3  G?�B�Y!dX   JJSr�3  G?�B�Y!duX   PRPr�3  j  �r�3  h h(h
c__builtin__
__main__
hNN}r�3  Ntr�3  Rr�3  �r�3  Rr�3  (h�G?�zoM�8X   VBPr�3  G?вB�YX   INr�3  G?вB�YX   NNr�3  G?�B�Y!dhMG?�B�Y!duX   NNSr�3  j�  �r�3  h h(h
c__builtin__
__main__
hNN}r�3  Ntr�3  Rr 4  �r4  Rr4  (h�G?�oM�7�X   INr4  G?��zoM�X   CDr4  G?�B�Y!dX   NNr4  G?�B�Y!dNG?�B�Y!dX   CCr4  G?�B�Y!dX   JJr4  G?�B�Y!dX   RBr4  G?�B�Y!dX   VBDr	4  G?�B�Y!dX   VBNr
4  G?�B�Y!dX   DTr4  G?�B�Y!dX   TOr4  G?�B�Y!dX   VBZr4  G?�B�Y!duX   NNr4  j�  �r4  h h(h
c__builtin__
__main__
hNN}r4  Ntr4  Rr4  �r4  Rr4  (X   RBr4  G?ѧ�a{�X   JJr4  G?�a{��h�G?��i�XGNG?���a{�X   INr4  G?���a{�X   VBNr4  G?���a{�X   NNSr4  G?���a{�X   NNr4  G?���a{�X   VBDr4  G?���a{�uj�  j4  �r4  h h(h
c__builtin__
__main__
hNN}r4  Ntr4  Rr4  �r 4  Rr!4  (X   VBNr"4  G?�Pה5�X   JJr#4  G?�򆼡�X   WPr$4  G?�򆼡�(h�G?�5�yC^X   VBZr%4  G?�5�yC^X   INr&4  G?�5�yC^X   VBr'4  G?�5�yC^X   VBGr(4  G?�򆼡�(X   VBPr)4  G?�ה5�yX   NNr*4  G?�򆼡�(X   VBDr+4  G?�����(lX   WRBr,4  G?�򆼡�(uX   DTr-4  j  �r.4  h h(h
c__builtin__
__main__
hNN}r/4  Ntr04  Rr14  �r24  Rr34  (X   NNSr44  G?�UUUUUUX   JJr54  G?�UUUUUUX   CDr64  G?�UUUUUUX   NNr74  G?�UUUUUUuX   WDTr84  j�  �r94  h h(h
c__builtin__
__main__
hNN}r:4  Ntr;4  Rr<4  �r=4  Rr>4  (X   RBr?4  G?�5�5�X   VBr@4  G?�@��@�X   DTrA4  G?�ЬЬX   JJrB4  G?�5�5�X   VBDrC4  G?�5�5�X   INrD4  G?�5�5�X   NNPrE4  G?�5�5�X   VBNrF4  G?�5�5�X   CCrG4  G?�5�5�uX   JJrH4  jW  �rI4  h h(h
c__builtin__
__main__
hNN}rJ4  NtrK4  RrL4  �rM4  RrN4  (X   NNrO4  G?�B�Y!X   JJrP4  G?ʶ�s��X   DTrQ4  G?���s��X   RBSrR4  G?���s��X   NNPrS4  G?�*K��a�X   NNSrT4  G?�B�Y!dX   NNPSrU4  G?�����X   TOrV4  G?�����X   VBZrW4  G?�����X   RBrX4  G?�����uX   VBGrY4  j�  �rZ4  h h(h
c__builtin__
__main__
hNN}r[4  Ntr\4  Rr]4  �r^4  Rr_4  (X   NNSr`4  G?��h�hX   INra4  G?�!�!�X   NNrb4  G?�����X   WPrc4  G?�!�!�X   VBGrd4  G?�����X   RBre4  G?�!�!�X   NNPrf4  G?��h�hX   CDrg4  G?���X   JJrh4  G?�!�!�X   VBNri4  G?���X   VBDrj4  G?��h�hX   DTrk4  G?��h�huX   MDrl4  j"  �rm4  h h(h
c__builtin__
__main__
hNN}rn4  Ntro4  Rrp4  �rq4  Rrr4  (X   VBGrs4  G?���k朐X   VBrt4  G?�NG�
�X   RBru4  G?�
�cp"X   WPrv4  G?�cp!���X   INrw4  G?�
�cp"X   JJrx4  G?���k朐X   MDry4  G?���k朐hMG?���k朐X   VBNrz4  G?���k朐X   VBPr{4  G?���k朐X   WDTr|4  G?���k朐uX   WRBr}4  hE�r~4  h h(h
c__builtin__
__main__
hNN}r4  Ntr�4  Rr�4  �r�4  Rr�4  (X   DTr�4  G?ϧ��~��X   JJr�4  G?��n[��X   NNr�4  G?�� HX   NNSr�4  G?�f��i�gX   VBZr�4  G?�@PX   PRPr�4  G?��0LX   NNPr�4  G?���|_�X   oovr�4  G?� @X   NNPSr�4  G?t@PX   VBr�4  G?� @X   JJSr�4  G?��p\X   RBr�4  G?���|X   RBSr�4  G?��0LX   VBNr�4  G?�� HX   CDr�4  G?|�pX   VBGr�4  G?�� HX   JJRr�4  G?� @X   VBDr�4  G?h�`X   ``r�4  G?` @uNh.�r�4  h h(h
c__builtin__
__main__
hNN}r�4  Ntr�4  Rr�4  �r�4  Rr�4  (X   NNSr�4  G?��e��l�X   VBPr�4  G?�
�B�P�X   INr�4  G?ȌF#��X   JJr�4  G?�M&�I��X   RBr�4  G?�
�B�P�X   NNr�4  G?����X   NNPr�4  G?����uj�  j�  �r�4  h h(h
c__builtin__
__main__
hNN}r�4  Ntr�4  Rr�4  �r�4  Rr�4  (X   JJr�4  G?�c�>pdX   PRPr�4  G?������X   WRBr�4  G?������X   RBr�4  G?������X   NNSr�4  G?������X   VBGr�4  G?�+��Q,X   DTr�4  G?�ډ]���X   NNr�4  G?������X   TOr�4  G?��Q+��X   INr�4  G?��Q+��X   PRP$r�4  G?������X   CCr�4  G?������X   VBNr�4  G?�81�8uX   WDTr�4  j1  �r�4  h h(h
c__builtin__
__main__
hNN}r�4  Ntr�4  Rr�4  �r�4  Rr�4  (X   NNSr�4  G?�X��Ƈ�X   JJr�4  G?�X��Ƈ�X   NNr�4  G?�Ƈ�4>�X   NNPr�4  G?�X��Ƈ�X   NNPSr�4  G?���/9X   CDr�4  G?�X��Ƈ�X   VBGr�4  G?���/9X   INr�4  G?���/9X   VBZr�4  G?���/9X   VBNr�4  G?���/9X   VBPr�4  G?���/9uX   NNSr�4  j�  �r�4  h h(h
c__builtin__
__main__
hNN}r�4  Ntr�4  Rr�4  �r�4  Rr�4  (X   NNr�4  G?���a{�h�G?�ܰ�=�	X   oovr�4  G?���a{�X   CCr�4  G?��i�XGhMG?���a{�X   NNPr�4  G?���a{�X   MDr�4  G?�{���aX   VBZr�4  G?���a{�X   VBDr�4  G?���a{�X   NNSr�4  G?���a|X   INr�4  G?���a{�X   VBPr�4  G?���a{�X   TOr�4  G?�{���aX   ``r�4  G?���a{�uNh/�r�4  h h(h
c__builtin__
__main__
hNN}r�4  Ntr�4  Rr�4  �r�4  Rr�4  (X   DTr�4  G?�Ǳ�{�X   NNr�4  G?��!�r�X   NNPr�4  G?����{��X   VBGr�4  G?�� HX   PRPr�4  G?��a�f�X   oovr�4  G?�$�2L�%X   VBNr�4  G?�� HX   JJr�4  G?�eYVU�eX   JJRr�4  G?h�`X   RBr�4  G?x�`X   NNPSr�4  G?h�`X   INr�4  G?h�`X   ``r�4  G?x�`X   CDr�4  G?h�`uX   VBNr�4  j�  �r�4  h h(h
c__builtin__
__main__
hNN}r�4  Ntr�4  Rr�4  �r�4  Rr�4  (X   NNr�4  G?�򆼡�(X   JJSr�4  G?�5�yC^X   JJr�4  G?�5�yC^X   NNSr�4  G?ǔ5�yCX   WPr�4  G?�򆼡�(X   CDr�4  G?�򆼡�(h�G?�򆼡�(uj�  j  �r�4  h h(h
c__builtin__
__main__
hNN}r�4  Ntr�4  Rr 5  �r5  Rr5  (X   VBr5  G?����8h#X   DTr5  G?���/��X   NNr5  G?���/��X   NNPr5  G?�[_u'X   NNPSr5  G?�[_u'uX   VBZr5  j�  �r	5  h h(h
c__builtin__
__main__
hNN}r
5  Ntr5  Rr5  �r5  Rr5  (X   VBr5  G?���ԇX   INr5  G?��+x�5X   TOr5  G?�MHs��X   VBZr5  G?�R�+x�X   VBNr5  G?����[�
h�G?·�R�X   JJr5  G?�&�9�V�X   CCr5  G?��+x�5"X   VBDr5  G?�R�+x�X   NNr5  G?�R�+x�X   WDTr5  G?����[�
X   VBPr5  G?��>��0MX   oovr5  G?|�+x�5"X   VBGr5  G?��+x�5"hMG?�&�9�V�X   NNSr5  G?�R�+x�X   RBr5  G?���[�	�X   DTr5  G?�&�9�V�X   MDr5  G?�R�+x�X   WRBr 5  G?�R�+x�X   POSr!5  G?��`����X   CDr"5  G?sR�+x�X   NNPr#5  G?sR�+x�ujN  j�  �r$5  h h(h
c__builtin__
__main__
hNN}r%5  Ntr&5  Rr'5  �r(5  Rr)5  (X   JJr*5  G?�zoM�8X   NNPr+5  G?��B�YX   VBGr,5  G?�B�Y!dh�G?�B�Y!dX   RBr-5  G?��B�YX   DTr.5  G?�B�Y!dX   PRPr/5  G?�B�Y!duhMj�"  �r05  h h(h
c__builtin__
__main__
hNN}r15  Ntr25  Rr35  �r45  Rr55  (X   INr65  G?�X   JJr75  G?�X   NNr85  G?�UUUUUUX   CCr95  G?ə�����X   NNPr:5  G?ə�����uX   ``r;5  j�%  �r<5  h h(h
c__builtin__
__main__
hNN}r=5  Ntr>5  Rr?5  �r@5  RrA5  (X   DTrB5  G?�UUUUUUX   PRPrC5  G?�UUUUUUX   INrD5  G?�      X   ''rE5  G?�UUUUUUX   TOrF5  G?�UUUUUUX   NNSrG5  G?�UUUUUUX   JJrH5  G?�      X   RBrI5  G?�UUUUUUX   VBNrJ5  G?�UUUUUUh�G?�UUUUUUuX   CDrK5  j`  �rL5  h h(h
c__builtin__
__main__
hNN}rM5  NtrN5  RrO5  �rP5  RrQ5  (h�G?�x���C�X   RBrR5  G?�`���ϚX   NNrS5  G?�x���C�X   JJrT5  G?��1��gX   TOrU5  G?�ԲN��X   NNSrV5  G?���@�hMG?�ԲN��X   NNPrW5  G?�`���ϚX   INrX5  G?�`���ϚX   VBNrY5  G?��1��gX   VBZrZ5  G?�`���ϚX   ``r[5  G?��1��gX   CCr\5  G?�2��tNG?�x���C�X   WRBr]5  G?��1��gX   WPr^5  G?�`���ϚX   CDr_5  G?�`���ϚX   JJSr`5  G?�`���ϚX   VBDra5  G?�`���ϚX   DTrb5  G?��1��gX   WDTrc5  G?�`���ϚX   PRPrd5  G?�`���ϚuX   WPre5  j\%  �rf5  h h(h
c__builtin__
__main__
hNN}rg5  Ntrh5  Rri5  �rj5  Rrk5  (X   NNrl5  G?�UUUUUUX   JJrm5  G?��8�9X   INrn5  G?�q�q�X   NNSro5  G?�UUUUUUuX   VBGrp5  hM�rq5  h h(h
c__builtin__
__main__
hNN}rr5  Ntrs5  Rrt5  �ru5  Rrv5  (X   VBGrw5  G?�zoM�8X   WRBrx5  G?��B�YX   WPry5  G?�zoM�8X   NNrz5  G?��zoM�X   INr{5  G?�B�Y!dX   CCr|5  G?��zoM�X   MDr}5  G?�B�Y!dX   VBZr~5  G?�B�Y!dX   DTr5  G?�B�Y!dX   CDr�5  G?�B�Y!duj)  j�  �r�5  h h(h
c__builtin__
__main__
hNN}r�5  Ntr�5  Rr�5  �r�5  Rr�5  (X   JJr�5  G?�      X   NNSr�5  G?�      X   CDr�5  G?�      X   NNr�5  G?�      h�G?�      X   NNPr�5  G?�      X   INr�5  G?�      uX   NNPSr�5  j  �r�5  h h(h
c__builtin__
__main__
hNN}r�5  Ntr�5  Rr�5  �r�5  Rr�5  (X   VBr�5  G?�      X   PRPr�5  G?�      X   DTr�5  G?�      X   NNr�5  G?�      X   RBr�5  G?�      X   TOr�5  G?�      ujt  j;&  �r�5  h h(h
c__builtin__
__main__
hNN}r�5  Ntr�5  Rr�5  �r�5  Rr�5  (X   JJr�5  G?��o��o�X   VBZr�5  G?�A�A�X   INr�5  G?�A�A�X   CDr�5  G?�UUUUUUX   NNSr�5  G?�A�A�X   VBNr�5  G?��;�;X   RBr�5  G?�i�i�X   DTr�5  G?�A�A�X   VBr�5  G?�A�A�X   VBPr�5  G?�A�A�uX   RPr�5  hM�r�5  h h(h
c__builtin__
__main__
hNN}r�5  Ntr�5  Rr�5  �r�5  Rr�5  (X   WPr�5  G?ə�����X   WRBr�5  G?�X   JJr�5  G?�X   MDr�5  G?�X   VBDr�5  G?�X   WDTr�5  G?�X   CCr�5  G?�uX   VBZr�5  j�
  �r�5  h h(h
c__builtin__
__main__
hNN}r�5  Ntr�5  Rr�5  �r�5  Rr�5  (X   VBr�5  G?�l�&ɲmX   DTr�5  G?�E�t]FX   RBr�5  G?�E�t]FX   NNPr�5  G?���|X   PRPr�5  G?�E�t]Fuj�  j+1  �r�5  h h(h
c__builtin__
__main__
hNN}r�5  Ntr�5  Rr�5  �r�5  Rr�5  (X   NNr�5  G?�2��s�X   INr�5  G?�lB:�I�X   NNPr�5  G?�+�_�j#h�G?��T{��VX   JJr�5  G?�Y�*tS6X   VBZr�5  G?k+�_�j#X   NNSr�5  G?�����$X   CDr�5  G?{+�_�j#X   CCr�5  G?��T{��VX   TOr�5  G?�`���ϚX   RBr�5  G?t`���ϚhMG?�+�_�j#X   ``r�5  G?k+�_�j#X   JJRr�5  G?t`���ϚX   WDTr�5  G?k+�_�j#X   VBr�5  G?��C��X   VBNr�5  G?�+�_�j#X   VBGr�5  G?k+�_�j#X   NNPSr�5  G?k+�_�j#X   DTr�5  G?k+�_�j#X   WPr�5  G?k+�_�j#X   POSr�5  G?k+�_�j#uX   VBZr�5  jR  �r�5  h h(h
c__builtin__
__main__
hNN}r�5  Ntr�5  Rr�5  �r�5  Rr�5  (X   INr�5  G?�dI囶X   JJr�5  G?�~�/�Q�X   VBPr�5  G?����X   DTr�5  G?�q|
���X   oovr�5  G?����Tt X   WPr�5  G?����X   RBr�5  G?����?WX   NNSr�5  G?����X   NNr�5  G?����Tt h�G?����X   VBZr�5  G?����X   CCr�5  G?����X   VBGr�5  G?����X   VBNr�5  G?����X   NNPr�5  G?����Tt X   CDr�5  G?����X   TOr�5  G?����X   ``r�5  G?����Tt X   PRPr�5  G?����hMG?����uX   oovr�5  jp&  �r�5  h h(h
c__builtin__
__main__
hNN}r�5  Ntr�5  Rr�5  �r�5  Rr�5  (X   VBPr�5  G?���HgoX   RBr�5  G?��֠R�[h�G?�&ɲl�'X   VBNr 6  G?��֠R�[hMG?���|X   CCr6  G?���|X   VBGr6  G?��֠R�[X   INr6  G?�&ɲl�'X   VBDr6  G?�q�q�X   JJr6  G?��֠R�[X   ''r6  G?��֠R�[X   NNSr6  G?��֠R�[X   TOr6  G?���|X   NNr	6  G?���|X   oovr
6  G?��֠R�[X   WRBr6  G?���|X   NNPr6  G?��֠R�[X   MDr6  G?���|uX   WPr6  j  �r6  h h(h
c__builtin__
__main__
hNN}r6  Ntr6  Rr6  �r6  Rr6  (X   NNSr6  G?���,�:h�G?�UUUUUUX   VBr6  G?��}�pX   DTr6  G?��tŝ1X   INr6  G?�򆼡�(X   VBNr6  G?�򆼡�(X   JJr6  G?�򆼡�(X   VBDr6  G?�򆼡�(X   VBPr6  G?�tŝ1gLX   NNr6  G?�򆼡�(X   PRPr6  G?��}�pX   CDr6  G?��}�pX   RBr 6  G?��}�pX   NNPr!6  G?�򆼡�(X   JJRr"6  G?��}�pX   RPr#6  G?�򆼡�(X   TOr$6  G?��}�pX   VBGr%6  G?��}�puX   VBr&6  ji  �r'6  h h(h
c__builtin__
__main__
hNN}r(6  Ntr)6  Rr*6  �r+6  Rr,6  (X   NNr-6  G?�I$�I$�X   VBGr.6  G?�a�a�X   NNPr/6  G?�I$�I$�X   JJSr06  G?�a�a�X   NNSr16  G?�y�y�X   JJr26  G?�a�a�X   INr36  G?�a�a�X   VBr46  G?�a�a�uX   WRBr56  hF�r66  h h(h
c__builtin__
__main__
hNN}r76  Ntr86  Rr96  �r:6  Rr;6  (X   DTr<6  G?ѧ�a{�X   NNPr=6  G?�/��JX   JJr>6  G?���lߢX   PRPr?6  G?��:ٿC�X   WRBr@6  G?w�L�x��X   JJSrA6  G?���a{�X   JJRrB6  G?��L�x��X   NNSrC6  G?�� ^)X   VBrD6  G?���a|X   VBNrE6  G?���a{�X   CDrF6  G?���a{�X   VBGrG6  G?���a{�X   NNrH6  G?���a|X   RBrI6  G?�lߡ���X   ``rJ6  G?w�L�x��X   NNPSrK6  G?���a{�X   PRP$rL6  G?w�L�x��h�G?w�L�x��uX   WDTrM6  j�  �rN6  h h(h
c__builtin__
__main__
hNN}rO6  NtrP6  RrQ6  �rR6  RrS6  (X   VBDrT6  G?�j%v�WjX   RBrU6  G?������X   VBPrV6  G?�#a�6#X   VBZrW6  G?����X   VBGrX6  G?������X   JJrY6  G?��Q+��X   NNPrZ6  G?���
h�X   CDr[6  G?���
h�X   VBNr\6  G?���
h�h�G?���
h�X   NNSr]6  G?������X   NNr^6  G?���
h�X   DTr_6  G?���
h�X   MDr`6  G?���
h�uX   RPra6  j�  �rb6  h h(h
c__builtin__
__main__
hNN}rc6  Ntrd6  Rre6  �rf6  Rrg6  (X   VBGrh6  G?�UUUUUUh�G?�      X   INri6  G?��q�rX   CDrj6  G?�q�q�X   TOrk6  G?�q�q�X   RBrl6  G?�q�q�X   VBPrm6  G?�q�q�X   JJrn6  G?�q�q�X   NNPro6  G?�q�q�uX   MDrp6  jP  �rq6  h h(h
c__builtin__
__main__
hNN}rr6  Ntrs6  Rrt6  �ru6  Rrv6  (h�G?�6�@�X   DTrw6  G?��V��X   PRP$rx6  G?��V��X   NNSry6  G?�Ի~2z�X   INrz6  G?�=K��'�X   NNr{6  G?�9��6X   VBr|6  G?� saZ$X   PRPr}6  G?��V��X   WPr~6  G?��V��X   VBGr6  G?��V��X   POSr�6  G?��V��X   RBr�6  G?��V��uX   MDr�6  j�  �r�6  h h(h
c__builtin__
__main__
hNN}r�6  Ntr�6  Rr�6  �r�6  Rr�6  (X   NNSr�6  G?�|��|X   NNr�6  G?�E�t]FX   NNPr�6  G?���|X   INr�6  G?�E�t]FX   NNPSr�6  G?���|X   JJr�6  G?�E�t]FX   DTr�6  G?���|X   VBGr�6  G?���|X   VBr�6  G?���|h�G?���|uX   JJSr�6  j  �r�6  h h(h
c__builtin__
__main__
hNN}r�6  Ntr�6  Rr�6  �r�6  Rr�6  (X   VBNr�6  G?�{���ahMG?�{���ah�G?���a|X   JJr�6  G?�ܰ�=�	X   VBr�6  G?���a{�X   INr�6  G?���a|X   VBGr�6  G?�{���aX   VBZr�6  G?���a{�X   VBPr�6  G?���a{�X   NNr�6  G?�{���aX   ''r�6  G?���a{�X   NNPr�6  G?�{���auX   NNPr�6  j	  �r�6  h h(h
c__builtin__
__main__
hNN}r�6  Ntr�6  Rr�6  �r�6  Rr�6  (X   CDr�6  G?��[���X   JJr�6  G?��[���X   DTr�6  G?�a2�aX   NNPr�6  G?��[���X   JJSr�6  G?��[���X   VBr�6  G?�*pA�*X   VBDr�6  G?�*pA�*X   NNr�6  G?�*pA�*X   VBGr�6  G?�m�ʜnh�G?�$�j��%X   INr�6  G?�a2�aX   CCr�6  G?��[���X   RBr�6  G?��[���X   VBNr�6  G?�m�ʜnNG?��[���X   NNSr�6  G?�m�ʜnX   WRBr�6  G?��[���uj	  j�6  �r�6  h h(h
c__builtin__
__main__
hNN}r�6  Ntr�6  Rr�6  �r�6  Rr�6  (X   INr�6  G?��w�GqX   NNPr�6  G?��_A}�X   CCr�6  G?��_A}�X   JJr�6  G?��_A}�X   NNr�6  G?��_A}�X   NNSr�6  G?��w�GqX   ''r�6  G?�_A}�X   JJSr�6  G?��_A}�X   ``r�6  G?��Gq�wX   oovr�6  G?��_A}�hMG?��_A}�uj�*  j2  �r�6  h h(h
c__builtin__
__main__
hNN}r�6  Ntr�6  Rr�6  �r�6  Rr�6  (h�G?��q�rX   NNSr�6  G?�UUUUUUX   INr�6  G?��q�rX   VBNr�6  G?��q�rX   VBr�6  G?�q�q�X   CCr�6  G?�q�q�X   DTr�6  G?�UUUUUUX   NNr�6  G?�UUUUUUX   VBPr�6  G?�UUUUUUuX   VBZr�6  j�!  �r�6  h h(h
c__builtin__
__main__
hNN}r�6  Ntr�6  Rr�6  �r�6  Rr�6  (X   NNSr�6  G?�B�Y!dX   RBr�6  G?�7��ޛ�X   JJr�6  G?�B�YX   VBNr�6  G?�B�Y!dX   VBr�6  G?�B�Y!dX   INr�6  G?��zoM�X   NNr�6  G?�B�Y!duX   ''r�6  j�  �r�6  h h(h
c__builtin__
__main__
hNN}r�6  Ntr�6  Rr�6  �r�6  Rr�6  (X   INr�6  G?��i�XGX   DTr�6  G?�ܰ�=�	X   WPr�6  G?���a{�X   RBr�6  G?�{���aX   VBNr�6  G?̰�=��X   WRBr�6  G?�{���aX   ``r�6  G?�{���aX   TOr�6  G?���a{�X   POSr�6  G?���a{�X   RPr�6  G?���a{�uj�  N�r�6  h h(h
c__builtin__
__main__
hNN}r�6  Ntr�6  Rr�6  �r�6  Rr�6  NG?�      sX   POSr�6  jZ  �r�6  h h(h
c__builtin__
__main__
hNN}r�6  Ntr�6  Rr 7  �r7  Rr7  (X   DTr7  G?�I$�I$�X   NNSr7  G?�m��m��X   CDr7  G?�m��m��X   NNPr7  G?�I$�I$�X   PRPr7  G?�I$�I$�h�G?�m��m��X   JJr7  G?�m��m��X   NNr	7  G?�m��m��X   oovr
7  G?�I$�I$�X   PRP$r7  G?�I$�I$�X   VBGr7  G?�m��m��X   WPr7  G?�I$�I$�uX   NNPSr7  hM�r7  h h(h
c__builtin__
__main__
hNN}r7  Ntr7  Rr7  �r7  Rr7  (X   NNPr7  G?�5�yC^X   WRBr7  G?�Pה5�X   WPr7  G?�򆼡�(X   NNPSr7  G?��5�yCX   VBDr7  G?�5�yC^X   INr7  G?�򆼡�(X   CCr7  G?�5�yC^X   WDTr7  G?�򆼡�(X   ''r7  G?�򆼡�(X   VBGr7  G?�򆼡�(X   DTr7  G?�5�yC^uX   RBr 7  j�  �r!7  h h(h
c__builtin__
__main__
hNN}r"7  Ntr#7  Rr$7  �r%7  Rr&7  (X   NNr'7  G?�X   INr(7  G?�/�b��0X   JJr)7  G?�N���OX   NNSr*7  G?�X   DTr+7  G?�N���OX   CDr,7  G?�N���OX   VBGr-7  G?�N���Oh�G?�X   VBNr.7  G?�N���OX   CCr/7  G?�z�G�{uX   TOr07  j  �r17  h h(h
c__builtin__
__main__
hNN}r27  Ntr37  Rr47  �r57  Rr67  (X   NNr77  G?�A�A�h�G?�m��m��X   INr87  G?��_�_X   VBDr97  G?�A�A�X   WPr:7  G?��_�_hMG?��_�_X   VBGr;7  G?�A�A�X   VBr<7  G?�A�A�uj�  j�/  �r=7  h h(h
c__builtin__
__main__
hNN}r>7  Ntr?7  Rr@7  �rA7  RrB7  (X   NNPrC7  G?��<��<�h�G?�m��m��X   VBrD7  G?�a�a�X   NNrE7  G?�a�a�X   NNSrF7  G?�a�a�X   CDrG7  G?�a�a�X   JJrH7  G?�a�a�X   oovrI7  G?�a�a�uj�  j�-  �rJ7  h h(h
c__builtin__
__main__
hNN}rK7  NtrL7  RrM7  �rN7  RrO7  (X   DTrP7  G?�333333X   VBrQ7  G?�������h�G?�X   WPrR7  G?�X   NNPrS7  G?�X   WDTrT7  G?�X   NNrU7  G?�X   RBrV7  G?�uX   VBNrW7  j�   �rX7  h h(h
c__builtin__
__main__
hNN}rY7  NtrZ7  Rr[7  �r\7  Rr]7  (X   VBNr^7  G?૰I���X   RBr_7  G?�v	2�:@X   MDr`7  G?����JX   oovra7  G?����JX   VBrb7  G?����JX   VBZrc7  G?���l֜\X   JJrd7  G?�TO�kNX   PRPre7  G?����JX   NNrf7  G?����JX   VBDrg7  G?��®�&SX   DTrh7  G?����JX   JJRri7  G?����JX   WPrj7  G?�e,t��7X   NNSrk7  G?�e,t��7X   VBGrl7  G?�e,t��7X   PRP$rm7  G?����JX   INrn7  G?�e,t��7X   VBPro7  G?�e,t��7X   WRBrp7  G?����JuX   JJrq7  jZ  �rr7  h h(h
c__builtin__
__main__
hNN}rs7  Ntrt7  Rru7  �rv7  Rrw7  (X   VBPrx7  G?�Y��Ig�X   NNSry7  G?��1�c�X   oovrz7  G?��`XX   INr{7  G?�2wH|��X   VBNr|7  G?�/��P��X   JJr}7  G?���f�\X   DTr~7  G?ν�z�X   JJSr7  G?���f�\X   NNr�7  G?�2wH|��X   JJRr�7  G?}\��ur�X   NNPr�7  G?�Y��Ig�X   VBGr�7  G?�\��ur�X   RBr�7  G?�\��ur�X   RPr�7  G?�\��ur�X   POSr�7  G?��`XX   PRPr�7  G?�Y��Ig�X   VBDr�7  G?��`XX   TOr�7  G?���f�\X   PRP$r�7  G?��`XX   CDr�7  G?}\��ur�X   MDr�7  G?}\��ur�X   VBr�7  G?��`XujZ  jx7  �r�7  h h(h
c__builtin__
__main__
hNN}r�7  Ntr�7  Rr�7  �r�7  Rr�7  (X   INr�7  G?�d�6M�eX   VBNr�7  G?�E�t]FX   JJr�7  G?���|X   WPr�7  G?���|X   NNSr�7  G?�E�t]FX   PRP$r�7  G?�E�t]FX   DTr�7  G?�E�t]FX   NNr�7  G?���|X   RBr�7  G?�E�t]FX   TOr�7  G?�E�t]FX   PRPr�7  G?���|uX   NNr�7  N�r�7  h h(h
c__builtin__
__main__
hNN}r�7  Ntr�7  Rr�7  �r�7  Rr�7  NG?�      sj�  j<&  �r�7  h h(h
c__builtin__
__main__
hNN}r�7  Ntr�7  Rr�7  �r�7  Rr�7  (X   NNSr�7  G?�TO�kNh�G?��®�&SX   INr�7  G?�v	2�:@X   WPr�7  G?�e,t��7X   PRPr�7  G?����JX   NNPr�7  G?����JX   VBGr�7  G?�e,t��7X   VBDr�7  G?����JX   TOr�7  G?�v	2�:@X   DTr�7  G?���D�f�X   NNr�7  G?��Ӌ<X   PRP$r�7  G?�e,t��7X   JJr�7  G?��Ӌ<X   VBNr�7  G?����JhMG?����JX   JJRr�7  G?�e,t��7X   RBr�7  G?����JX   WDTr�7  G?����JX   VBPr�7  G?�e,t��7X   CDr�7  G?����JX   VBr�7  G?����JuX   CDr�7  N�r�7  h h(h
c__builtin__
__main__
hNN}r�7  Ntr�7  Rr�7  �r�7  Rr�7  NG?�      sj�   j�,  �r�7  h h(h
c__builtin__
__main__
hNN}r�7  Ntr�7  Rr�7  �r�7  Rr�7  (X   VBr�7  G?��I�A�X   JJr�7  G?�[_u'X   NNPr�7  G?���/��h�G?�_u'WX   WRBr�7  G?���/��X   WPr�7  G?�[_u'X   DTr�7  G?�_u'WX   CDr�7  G?�[_u'X   NNSr�7  G?�[_u'X   INr�7  G?���/��X   RBr�7  G?�[_u'uX   NNPSr�7  j3  �r�7  h h(h
c__builtin__
__main__
hNN}r�7  Ntr�7  Rr�7  �r�7  Rr�7  (X   RPr�7  G?�UUUUUUX   INr�7  G?�UUUUUUX   NNPr�7  G?�������X   NNr�7  G?�UUUUUUh�G?�������X   DTr�7  G?ª�����X   TOr�7  G?ª�����X   POSr�7  G?�UUUUUUX   NNSr�7  G?�UUUUUUX   JJr�7  G?�UUUUUUX   PRP$r�7  G?�UUUUUUX   WPr�7  G?�UUUUUUuX   VBPr�7  j�  �r�7  h h(h
c__builtin__
__main__
hNN}r�7  Ntr�7  Rr�7  �r�7  Rr�7  (X   JJr�7  G?�>�>�X   DTr�7  G?�>�>�X   NNPr�7  G?�>�>�X   INr�7  G?�&=�&=�h�G?���X   NNr�7  G?�N�N�X   VBNr�7  G?��$�$X   PRP$r�7  G?�~h~hX   RPr�7  G?�~h~hX   NNSr�7  G?�֒�֒�X   POSr�7  G?�����X   TOr�7  G?�~h~hX   WPr�7  G?�~h~hX   CCr�7  G?�~h~hX   JJRr�7  G?�����X   RBr�7  G?��$�$X   oovr�7  G?�>�>�X   WRBr�7  G?�����X   PRPr 8  G?�����X   VBGr8  G?�����NG?�����X   VBr8  G?�����uX   NNPSr8  j3  �r8  h h(h
c__builtin__
__main__
hNN}r8  Ntr8  Rr8  �r8  Rr	8  (X   DTr
8  G?�m��m��h�G?ĒI$�I%X   INr8  G?�      X   TOr8  G?�m��m��X   JJr8  G?��m��m�X   NNSr8  G?�m��m��X   NNPr8  G?�I$�I$�X   PRPr8  G?�m��m��X   NNr8  G?��m��m�X   PRP$r8  G?�      X   VBNr8  G?�      X   WRBr8  G?�I$�I$�X   VBGr8  G?�I$�I$�X   RBr8  G?�I$�I$�X   NNPSr8  G?�I$�I$�X   RPr8  G?�I$�I$�X   JJRr8  G?�I$�I$�X   WDTr8  G?�I$�I$�X   VBZr8  G?�I$�I$�X   oovr8  G?�I$�I$�uX   RPr8  j  �r8  h h(h
c__builtin__
__main__
hNN}r8  Ntr 8  Rr!8  �r"8  Rr#8  (h�G?͉؝�؞X   INr$8  G?؝�؝��X   TOr%8  G?��؝�؞X   NNSr&8  G?��;�;X   VBPr'8  G?��;�;X   CCr(8  G?��;�;X   DTr)8  G?��;�;X   VBGr*8  G?��;�;X   VBr+8  G?��;�;X   VBDr,8  G?��؝�؞uX   DTr-8  j�  �r.8  h h(h
c__builtin__
__main__
hNN}r/8  Ntr08  Rr18  �r28  Rr38  (X   VBPr48  G?�'�n�i�X   INr58  G?����h�G?�_���\X   VBDr68  G?����Tt X   RBr78  G?����X   MDr88  G?����X   VBZr98  G?����Tt X   NNr:8  G?�yf톙X   JJr;8  G?����Tt X   ''r<8  G?����uX   NNPSr=8  j  �r>8  h h(h
c__builtin__
__main__
hNN}r?8  Ntr@8  RrA8  �rB8  RrC8  (X   DTrD8  G?��w�GqX   WDTrE8  G?��_A}�X   NNPrF8  G?��_A}�X   INrG8  G?��SYMe6X   PRP$rH8  G?��_A}�X   VBNrI8  G?��_A}�X   RBrJ8  G?��Gq�wX   WRBrK8  G?��_A}�X   WPrL8  G?��_A}�X   JJrM8  G?��Gq�wX   NNrN8  G?��_A}�X   PRPrO8  G?��_A}�uX   NNPSrP8  j  �rQ8  h h(h
c__builtin__
__main__
hNN}rR8  NtrS8  RrT8  �rU8  RrV8  (h�G?��V��X   RPrW8  G?��V��X   VBNrX8  G?��@�´HX   NNrY8  G?��V��X   INrZ8  G?�$l+D�X   DTr[8  G?��V��X   TOr\8  G?�6�@�X   VBGr]8  G?��V��X   oovr^8  G?��V��uX   VBZr_8  jE8  �r`8  h h(h
c__builtin__
__main__
hNN}ra8  Ntrb8  Rrc8  �rd8  Rre8  (X   NNrf8  G?ׂ����X   INrg8  G?�X��ƈX   VBGrh8  G?���/9X   NNSri8  G?�X��Ƈ�X   NNPrj8  G?���/9X   CDrk8  G?���/9X   VBDrl8  G?���/9X   VBPrm8  G?�X��ƈX   JJrn8  G?���/9X   MDro8  G?���/9X   VBrp8  G?���/9X   VBZrq8  G?���/9uX   DTrr8  j�  �rs8  h h(h
c__builtin__
__main__
hNN}rt8  Ntru8  Rrv8  �rw8  Rrx8  (X   DTry8  G?�t]E�tX   VBZrz8  G?��A)��X   INr{8  G?�E�t]FX   JJr|8  G?��A)��h�G?�Jy��JX   NNr}8  G?�Jy��JX   WPr~8  G?��A)��X   NNSr8  G?��A)��X   VBNr�8  G?��A)��X   RBr�8  G?��A)��X   ``r�8  G?�E�t]FuX   JJr�8  j�  �r�8  h h(h
c__builtin__
__main__
hNN}r�8  Ntr�8  Rr�8  �r�8  Rr�8  (X   VBDr�8  G?�3�* hX   INr�8  G?�* g�:TX   NNr�8  G?�쎕3�h�G?�3�* hX   JJr�8  G?�쎕3�X   NNSr�8  G?�쎕3�X   DTr�8  G?�쎕3�X   VBPr�8  G?�쎕3�hMG?�쎕3�X   VBZr�8  G?�쎕3�uj  j�"  �r�8  h h(h
c__builtin__
__main__
hNN}r�8  Ntr�8  Rr�8  �r�8  Rr�8  (X   NNPr�8  G?�      X   CDr�8  G?�      X   NNr�8  G?�      X   JJr�8  G?�      uX   NNPSr�8  j	  �r�8  h h(h
c__builtin__
__main__
hNN}r�8  Ntr�8  Rr�8  �r�8  Rr�8  (X   JJr�8  G?��m��m�X   NNSr�8  G?�I$�I$�X   NNPr�8  G?�I$�I$�X   NNr�8  G?�m��m��X   JJSr�8  G?�m��m��h�G?�m��m��X   NNPSr�8  G?�m��m��uX   NNPSr�8  j
  �r�8  h h(h
c__builtin__
__main__
hNN}r�8  Ntr�8  Rr�8  �r�8  Rr�8  (X   VBr�8  G?��ͣ�X   VBPr�8  G?��qO��;h�G?��qO��;X   TOr�8  G?��ͣ��X   INr�8  G?��qO��;X   RBr�8  G?��qO��;X   JJr�8  G?�.)��GXX   VBNr�8  G?�.)��GXX   VBDr�8  G?�.)��GXuX   INr�8  j=  �r�8  h h(h
c__builtin__
__main__
hNN}r�8  Ntr�8  Rr�8  �r�8  Rr�8  (X   NNr�8  G?�[_u'X   VBPr�8  G?�[_u'h�G?�z�$(X   VBGr�8  G?�[_u'X   VBNr�8  G?�?�o^�X   VBDr�8  G?�ѷ�rCX   WPr�8  G?�$(F޼X   INr�8  G?�_u'WX   DTr�8  G?�$(F޼X   POSr�8  G?�[_u'X   TOr�8  G?�$(F޼X   NNPr�8  G?�$(F޼X   CCr�8  G?�ѷ�rCX   JJr�8  G?�[_u'hMG?�$(F޼X   ''r�8  G?�[_u'X   NNSr�8  G?�[_u'X   CDr�8  G?�$(F޼X   VBr�8  G?��2��kX   WRBr�8  G?�$(F޼X   VBZr�8  G?�$(F޼X   RBr�8  G?�[_u'uX   JJr�8  j\  �r�8  h h(h
c__builtin__
__main__
hNN}r�8  Ntr�8  Rr�8  �r�8  Rr�8  (X   VBDr�8  G?��� OX   VBNr�8  G?�9&\a�h�G?�Z�>�E�X   VBPr�8  G?��])~X   INr�8  G?�#:�1R4X   NNSr�8  G?��/�^�X   NNPr�8  G?���M�,�X   NNr�8  G?�|z �w�X   WPr�8  G?���M�,�X   RBr�8  G?��/�^�X   CCr�8  G?���M�,�X   VBr�8  G?���M�,�X   JJr�8  G?���M�,�X   ''r�8  G?�O��hMG?�O��X   oovr�8  G?yO��X   TOr�8  G?�O��X   VBGr�8  G?���M�,�X   NNPSr�8  G?yO��X   VBZr�8  G?�O��X   DTr�8  G?���M�,�X   MDr�8  G?���M�,�X   POSr�8  G?���M�,�X   ``r�8  G?�P�ց�
uX   JJr�8  j�  �r�8  h h(h
c__builtin__
__main__
hNN}r�8  Ntr�8  Rr�8  �r�8  Rr�8  (X   RBr�8  G?�      X   JJr�8  G?⪪����X   NNr�8  G?�      X   VBGr�8  G?�UUUUUUX   NNPSr�8  G?�UUUUUUX   VBNr�8  G?�      X   NNSr�8  G?�UUUUUUX   NNPr�8  G?�UUUUUUuX   VBZr�8  jV  �r 9  h h(h
c__builtin__
__main__
hNN}r9  Ntr9  Rr9  �r9  Rr9  (X   JJSr9  G?�ЬЬX   TOr9  G?�X   JJr9  G?�ЬЬX   DTr	9  G?�oݔoݔX   INr
9  G?�ЬЬh�G?��:�:X   VBGr9  G?�ЬЬX   NNPr9  G?�5�5�X   NNSr9  G?��:�:X   oovr9  G?�5�5�X   RBr9  G?��:�:X   WPr9  G?��:�:X   CDr9  G?�5�5�X   PRP$r9  G?�5�5�X   NNr9  G?�5�5�X   JJRr9  G?�5�5�ujV  j9  �r9  h h(h
c__builtin__
__main__
hNN}r9  Ntr9  Rr9  �r9  Rr9  (X   INr9  G?�333333X   NNr9  G?�X   NNSr9  G?�X   JJr9  G?�uj�8  j$  �r9  h h(h
c__builtin__
__main__
hNN}r 9  Ntr!9  Rr"9  �r#9  Rr$9  (X   JJr%9  G?؝�؝��X   RBr&9  G?��o��o�X   INr'9  G?�A�A�h�G?�A�A�X   VBNr(9  G?�A�A�X   VBPr)9  G?�A�A�X   NNr*9  G?�A�A�uX   NNPr+9  j	  �r,9  h h(h
c__builtin__
__main__
hNN}r-9  Ntr.9  Rr/9  �r09  Rr19  (X   RBr29  G?�UUUUUUX   JJr39  G?�&ɲl�'X   VBr49  G?���|X   VBNr59  G?�E�t]FX   VBDr69  G?�E�t]FuhMj�  �r79  h h(h
c__builtin__
__main__
hNN}r89  Ntr99  Rr:9  �r;9  Rr<9  (X   RBr=9  G?�c�qF:�X   NNSr>9  G?�/�A��4X   CCr?9  G?���!�xhMG?���!�xX   VBNr@9  G?�A��40X   NNPrA9  G?���!�xX   VBPrB9  G?���!�xX   WPrC9  G?�/�A��4X   INrD9  G?���ajzVX   DTrE9  G?Ņ��XZ�X   NNrF9  G?���!�xX   JJRrG9  G?���!�xX   VBZrH9  G?���!�xX   PRPrI9  G?�/�A��4X   CDrJ9  G?���!�xX   JJrK9  G?�/�A��4X   RPrL9  G?���!�xX   PRP$rM9  G?�/�A��4X   VBrN9  G?���!�xX   WRBrO9  G?�/�A��4X   VBDrP9  G?���!�xX   RBSrQ9  G?�/�A��4X   VBGrR9  G?���!�xX   JJSrS9  G?���!�xuX   MDrT9  j  �rU9  h h(h
c__builtin__
__main__
hNN}rV9  NtrW9  RrX9  �rY9  RrZ9  (X   NNPr[9  G?�&��h�'X   VBr\9  G?ֵ�kZֶX   POSr]9  G?ĥ)JR��X   CCr^9  G?��!B�X   NNSr_9  G?��`XX   RBr`9  G?��!B�h�G?��`XX   NNra9  G?���n�X   VBDrb9  G?��`XuX   RPrc9  j�  �rd9  h h(h
c__builtin__
__main__
hNN}re9  Ntrf9  Rrg9  �rh9  Rri9  (X   NNSrj9  G?θQ��X   VBrk9  G?�z�G�{X   TOrl9  G?�z�G�{X   CCrm9  G?��Q��X   NNrn9  G?�333333X   JJro9  G?���Q�X   NNPrp9  G?�������X   INrq9  G?�z�G�{uX   VBPrr9  j�  �rs9  h h(h
c__builtin__
__main__
hNN}rt9  Ntru9  Rrv9  �rw9  Rrx9  (h�G?������X   VBry9  G?�j%v�WjX   VBNrz9  G?�81�8X   RBr{9  G?�81�8X   VBGr|9  G?��Q+��X   INr}9  G?������X   VBDr~9  G?��Q+��X   CDr9  G?������X   DTr�9  G?������uX   RPr�9  j�  �r�9  h h(h
c__builtin__
__main__
hNN}r�9  Ntr�9  Rr�9  �r�9  Rr�9  (X   NNr�9  G?�E�t]h�G?�t]E�tX   RBr�9  G?�E�t]FX   VBGr�9  G?�E�t]FX   INr�9  G?�E�t]FX   NNSr�9  G?�t]E�tX   JJr�9  G?�E�t]FX   NNPr�9  G?�E�t]FX   PRPr�9  G?�E�t]FX   VBZr�9  G?�t]E�tuj=.  j0  �r�9  h h(h
c__builtin__
__main__
hNN}r�9  Ntr�9  Rr�9  �r�9  Rr�9  (X   CDr�9  G?��u�u h�G?��p�pX   VBNr�9  G?��p�pX   NNr�9  G?��k�kX   INr�9  G?�l�l�X   oovr�9  G?�PPPPPPX   NNPr�9  G?�X   RBr�9  G?��p�pX   VBDr�9  G?�X   NNSr�9  G?��p�pX   JJSr�9  G?��p�pX   JJr�9  G?�X   VBZr�9  G?��p�phMG?��p�pX   CCr�9  G?��p�pNG?�X   DTr�9  G?��p�puhMju  �r�9  h h(h
c__builtin__
__main__
hNN}r�9  Ntr�9  Rr�9  �r�9  Rr�9  (X   WPr�9  G?�m��m��X   NNSr�9  G?�A�A�X   VBr�9  G?�I$�I$�X   PRP$r�9  G?�A�A�X   RBr�9  G?��_�_X   WRBr�9  G?��_�_uX   WPr�9  j�  �r�9  h h(h
c__builtin__
__main__
hNN}r�9  Ntr�9  Rr�9  �r�9  Rr�9  (X   NNr�9  G?�UUUUUUX   VBZr�9  G?�UUUUUUX   JJr�9  G?�UUUUUUh�G?�UUUUUUX   INr�9  G?�UUUUUUuX   WRBr�9  j  �r�9  h h(h
c__builtin__
__main__
hNN}r�9  Ntr�9  Rr�9  �r�9  Rr�9  (X   NNPr�9  G?�X   VBPr�9  G?�X   NNSr�9  G?�333333X   NNr�9  G?�������X   VBZr�9  G?�X   JJr�9  G?�X   CCr�9  G?�X   VBDr�9  G?�X   INr�9  G?�uX   WPr�9  jq  �r�9  h h(h
c__builtin__
__main__
hNN}r�9  Ntr�9  Rr�9  �r�9  Rr�9  (X   NNPr�9  G?�����/hX   INr�9  G?�q�q�X   NNr�9  G?ք��/hLX   VBDr�9  G?��%�	{BX   VBPr�9  G?�����/hX   VBGr�9  G?�����/hX   JJr�9  G?�����/hX   DTr�9  G?�q�q�X   RBr�9  G?�����/hX   JJRr�9  G?�����/hX   RBSr�9  G?�����/hX   VBZr�9  G?�����/huh�j�  �r�9  h h(h
c__builtin__
__main__
hNN}r�9  Ntr�9  Rr�9  �r�9  Rr�9  (X   VBPr�9  G?�      X   VBZr�9  G?�UUUUUUX   VBDr�9  G?�      X   NNr�9  G?�UUUUUUuX   JJSr�9  hM�r�9  h h(h
c__builtin__
__main__
hNN}r�9  Ntr�9  Rr�9  �r�9  Rr�9  (X   JJSr�9  G?�UUUUUUX   INr�9  G?�      X   MDr�9  G?�UUUUUUX   RBSr�9  G?�      X   NNr�9  G?�UUUUUUuhMj�9  �r�9  h h(h
c__builtin__
__main__
hNN}r�9  Ntr�9  Rr�9  �r�9  Rr�9  (X   NNr�9  G?�t]E�tX   NNSr�9  G?�t]E�tX   PRPr�9  G?�E�t]FX   JJr�9  G?�t]E�tuj�  j�8  �r�9  h h(h
c__builtin__
__main__
hNN}r :  Ntr:  Rr:  �r:  Rr:  (X   NNSr:  G?���SF�X   VBNr:  G?���:�7�X   VBDr:  G?���ː��X   INr:  G?Ǆ�b��>X   DTr	:  G?�Yr��SX   NNPr
:  G?�F�V]X   PRP$r:  G?��P1YrX   NNr:  G?��!�~u4X   TOr:  G?��SF�h�G?�7��b��X   RBr:  G?��P1YrX   RPr:  G?���k�X   JJr:  G?�1Yr��X   oovr:  G?���ː��X   CDr:  G?x��k�X   WPr:  G?x��k�X   WRBr:  G?���ː��X   PRPr:  G?���SF�X   VBGr:  G?���k�X   WDTr:  G?x��k�uX   VBPr:  j
  �r:  h h(h
c__builtin__
__main__
hNN}r:  Ntr:  Rr:  �r:  Rr:  (h�G?�X   VBDr:  G?ə�����X   VBPr :  G?�������X   VBr!:  G?�X   INr":  G?�X   NNr#:  G?�X   MDr$:  G?�������X   NNSr%:  G?�X   VBZr&:  G?ə�����uj
  h��r':  h h(h
c__builtin__
__main__
hNN}r(:  Ntr):  Rr*:  �r+:  Rr,:  NG?�      sX   NNSr-:  j#  �r.:  h h(h
c__builtin__
__main__
hNN}r/:  Ntr0:  Rr1:  �r2:  Rr3:  (X   INr4:  G?θQ��X   NNr5:  G?ə�����X   CCr6:  G?�z�G�{h�G?�z�G�{X   NNSr7:  G?�z�G�{X   RBr8:  G?�z�G�{X   WPr9:  G?�z�G�{X   PRPr::  G?�z�G�{uX   VBPr;:  j  �r<:  h h(h
c__builtin__
__main__
hNN}r=:  Ntr>:  Rr?:  �r@:  RrA:  (X   JJrB:  G?�m��m��X   VBNrC:  G?�I$�I$�X   VBrD:  G?ĒI$�I%X   RBrE:  G?�I$�I$�X   NNSrF:  G?�$�I$�IX   NNPrG:  G?�m��m��X   NNrH:  G?�I$�I$�X   JJRrI:  G?�I$�I$�uX   CDrJ:  jS  �rK:  h h(h
c__builtin__
__main__
hNN}rL:  NtrM:  RrN:  �rO:  RrP:  (X   VBNrQ:  G?�X   NNSrR:  G?�X   DTrS:  G?�X   JJRrT:  G?�X   PRP$rU:  G?�X   INrV:  G?�X   WPrW:  G?�X   JJrX:  G?�X   TOrY:  G?�X   WRBrZ:  G?�h�G?�X   RBr[:  G?�X   NNPr\:  G?�X   NNr]:  G?�uX   MDr^:  j   �r_:  h h(h
c__builtin__
__main__
hNN}r`:  Ntra:  Rrb:  �rc:  Rrd:  (X   VBre:  G?�؝�؞X   POSrf:  G?��;�;X   NNrg:  G?�;�;�X   ``rh:  G?��;�;X   JJRri:  G?��;�;X   NNSrj:  G?��؝�؞X   JJrk:  G?��;�;X   RBrl:  G?��;�;X   VBZrm:  G?��;�;X   INrn:  G?��;�;uX   CCro:  j�  �rp:  h h(h
c__builtin__
__main__
hNN}rq:  Ntrr:  Rrs:  �rt:  Rru:  (h�G?�UUUUUUX   VBZrv:  G?ə�����X   TOrw:  G?�X   RBrx:  G?�X   VBDry:  G?�X   NNrz:  G?�NG?�X   VBPr{:  G?�UUUUUUX   MDr|:  G?�uX   RBSr}:  jC:  �r~:  h h(h
c__builtin__
__main__
hNN}r:  Ntr�:  Rr�:  �r�:  Rr�:  (X   INr�:  G?�v'bv'bX   TOr�:  G?��؝�؞h�G?ȝ�؝��X   WRBr�:  G?��؝�؞uj�  jh8  �r�:  h h(h
c__builtin__
__main__
hNN}r�:  Ntr�:  Rr�:  �r�:  Rr�:  (X   NNSr�:  G?�UUUUUUX   NNr�:  G?�UUUUUUX   NNPr�:  G?�UUUUUUh�G?�UUUUUUuX   DTr�:  j�  �r�:  h h(h
c__builtin__
__main__
hNN}r�:  Ntr�:  Rr�:  �r�:  Rr�:  (X   NNr�:  G?�I$�I$�X   VBDr�:  G?�I$�I$�X   TOr�:  G?�I$�I$�X   VBPr�:  G?�I$�I$�X   VBZr�:  G?�I$�I$�X   DTr�:  G?�I$�I$�uNh0�r�:  h h(h
c__builtin__
__main__
hNN}r�:  Ntr�:  Rr�:  �r�:  Rr�:  (X   DTr�:  G?�UUUUUUX   NNSr�:  G?�H+�d�X   PRPr�:  G?��l�lX   RBr�:  G?��l�lX   RBSr�:  G?��l�lX   JJr�:  G?���j1M�X   PRP$r�:  G?�W:��tX   oovr�:  G?�����/hX   JJRr�:  G?�W:��tX   VBNr�:  G?��l�lX   ``r�:  G?��l�luX   VBr�:  h��r�:  h h(h
c__builtin__
__main__
hNN}r�:  Ntr�:  Rr�:  �r�:  Rr�:  (X   VBr�:  G?��/���X   DTr�:  G?��_A}�X   RBr�:  G?��Gq�wuX   VBZr�:  j�!  �r�:  h h(h
c__builtin__
__main__
hNN}r�:  Ntr�:  Rr�:  �r�:  Rr�:  (X   VBZr�:  G?�      X   DTr�:  G?�򆼡�(X   NNSr�:  G?ǔ5�yCX   JJRr�:  G?�򆼡�(X   VBr�:  G?�򆼡�(X   NNr�:  G?�򆼡�(X   RBr�:  G?�򆼡�(uX   NNSr�:  j�  �r�:  h h(h
c__builtin__
__main__
hNN}r�:  Ntr�:  Rr�:  �r�:  Rr�:  (X   INr�:  G?��"�TX   CCr�:  G?�k݀�fX   JJr�:  G?����"X   DTr�:  G?���n�tX   NNr�:  G?�'�y�8IX   ``r�:  G?���n�tX   RBr�:  G?�'�y�8IX   VBZr�:  G?���n�tX   NNPSr�:  G?���n�tX   NNSr�:  G?�Ɉ+�WX   WPr�:  G?�Ɉ+�WX   VBr�:  G?���n�thMG?���n�th�G?���n�tX   VBNr�:  G?���n�tX   ''r�:  G?���n�tX   VBGr�:  G?���n�tX   TOr�:  G?���n�tX   VBPr�:  G?���n�tX   NNPr�:  G?�Ɉ+�WX   CDr�:  G?���n�tX   VBDr�:  G?���n�tNG?���n�tuX   PRPr�:  j�  �r�:  h h(h
c__builtin__
__main__
hNN}r�:  Ntr�:  Rr�:  �r�:  Rr�:  (X   DTr�:  G?�d�6M�eX   JJr�:  G?���|X   VBNr�:  G?���|X   NNPr�:  G?���|h�G?���|X   VBr�:  G?���|X   INr�:  G?���|X   VBZr�:  G?���|X   WRBr�:  G?���|X   RBr�:  G?���|uh�h��r�:  h h(h
c__builtin__
__main__
hNN}r�:  Ntr�:  Rr�:  �r�:  Rr�:  (NG?��h�2\X   INr�:  G?��qO��;uhMj�  �r�:  h h(h
c__builtin__
__main__
hNN}r�:  Ntr�:  Rr�:  �r�:  Rr�:  (X   NNr�:  G?�UUUUUUX   NNSr�:  G?�q�q�X   JJr ;  G?�q�q�uX   JJSr;  j  �r;  h h(h
c__builtin__
__main__
hNN}r;  Ntr;  Rr;  �r;  Rr;  (X   MDr;  G?�      X   VBPr	;  G?�      X   NNSr
;  G?�      h�G?�      uX   WRBr;  j�4  �r;  h h(h
c__builtin__
__main__
hNN}r;  Ntr;  Rr;  �r;  Rr;  (X   PRPr;  G?�I$�I$�X   DTr;  G?�m��m��X   RBr;  G?�I$�I$�uj  j�:  �r;  h h(h
c__builtin__
__main__
hNN}r;  Ntr;  Rr;  �r;  Rr;  (X   oovr;  G?݉؝�؞X   JJRr;  G?ȝ�؝��X   DTr;  G?�A�A�X   VBGr;  G?�A�A�X   NNPr;  G?�A�A�X   NNr ;  G?�A�A�hMG?�A�A�X   VBr!;  G?�A�A�X   VBNr";  G?�A�A�X   CDr#;  G?�A�A�X   JJr$;  G?�A�A�X   RBr%;  G?�A�A�X   CCr&;  G?��;�;X   PRPr';  G?�A�A�uNh1�r(;  h h(h
c__builtin__
__main__
hNN}r);  Ntr*;  Rr+;  �r,;  Rr-;  (X   INr.;  G?�UUUUUUX   JJr/;  G?�q�q�X   NNr0;  G?�q�q�X   NNSr1;  G?�q�q�uX   PRP$r2;  j�  �r3;  h h(h
c__builtin__
__main__
hNN}r4;  Ntr5;  Rr6;  �r7;  Rr8;  X   JJr9;  G?�      sX   POSr:;  jR5  �r;;  h h(h
c__builtin__
__main__
hNN}r<;  Ntr=;  Rr>;  �r?;  Rr@;  (X   VBNrA;  G?�ֵ�kZ�X   VBPrB;  G?��1�c�X   JJrC;  G?��1�c�X   VBGrD;  G?��!B�X   VBrE;  G?��1�c�X   NNPrF;  G?��!B�uh�j�  �rG;  h h(h
c__builtin__
__main__
hNN}rH;  NtrI;  RrJ;  �rK;  RrL;  (X   CDrM;  G?�t]E�tX   NNPrN;  G?�]E�t]X   NNrO;  G?�t]E�tX   VBPrP;  G?�E�t]FX   POSrQ;  G?�.���/hMG?�E�t]Fh�G?�t]E�tX   CCrR;  G?�E�t]FX   VBDrS;  G?�t]E�tX   VBrT;  G?�t]E�tX   JJrU;  G?�E�t]FX   DTrV;  G?�t]E�tX   VBGrW;  G?�E�t]FX   RBrX;  G?�E�t]FX   VBNrY;  G?�E�t]FX   VBZrZ;  G?�E�t]FX   INr[;  G?�E�t]FuX   JJr\;  j�  �r];  h h(h
c__builtin__
__main__
hNN}r^;  Ntr_;  Rr`;  �ra;  Rrb;  (X   DTrc;  G?ñ;�;X   INrd;  G?͉؝�؞h�G?ӱ;�;X   POSre;  G?ñ;�;X   NNPrf;  G?ñ;�;uX   POSrg;  j[  �rh;  h h(h
c__builtin__
__main__
hNN}ri;  Ntrj;  Rrk;  �rl;  Rrm;  (X   NNPrn;  G?�[�[�X   NNro;  G?�X   JJrp;  G?�X   VBZrq;  G?��l�lX   NNSrr;  G?�X   CCrs;  G?��l�luj�,  j�#  �rt;  h h(h
c__builtin__
__main__
hNN}ru;  Ntrv;  Rrw;  �rx;  Rry;  (X   RBrz;  G?�(�\)X   VBr{;  G?�
=p��
X   DTr|;  G?�z�G�{X   PRPr};  G?��Q��uX   ``r~;  j�  �r;  h h(h
c__builtin__
__main__
hNN}r�;  Ntr�;  Rr�;  �r�;  Rr�;  (X   CDr�;  G?����� X   VBGr�;  G?��z�zX   DTr�;  G?��z�zX   JJr�;  G?ˑ���X   ''r�;  G?ǡz�zX   RBr�;  G?��;�;X   PRPr�;  G?����� X   VBNr�;  G?��z�zhMG?��z�zX   INr�;  G?��z�zX   TOr�;  G?����� X   NNr�;  G?����� h�G?��z�zX   PRP$r�;  G?����� X   ``r�;  G?����� X   VBZr�;  G?����� uj�;  jf2  �r�;  h h(h
c__builtin__
__main__
hNN}r�;  Ntr�;  Rr�;  �r�;  Rr�;  (h�G?ə�����NG?�������hMG?�������X   VBZr�;  G?�������X   NNr�;  G?�333333X   VBDr�;  G?�333333X   VBNr�;  G?�������X   VBr�;  G?�333333X   NNSr�;  G?�������uh�jl3  �r�;  h h(h
c__builtin__
__main__
hNN}r�;  Ntr�;  Rr�;  �r�;  Rr�;  (X   JJr�;  G?ə�����X   RBSr�;  G?�X   NNPr�;  G?ə�����X   NNr�;  G?�������uX   PRP$r�;  j�  �r�;  h h(h
c__builtin__
__main__
hNN}r�;  Ntr�;  Rr�;  �r�;  Rr�;  (X   RBSr�;  G?�a�a�X   NNr�;  G?�y�y�X   JJSr�;  G?�a�a�X   NNPr�;  G?�a�a�X   JJr�;  G?�I$�I$�X   INr�;  G?�I$�I$�X   VBGr�;  G?�a�a�uj�  j�;  �r�;  h h(h
c__builtin__
__main__
hNN}r�;  Ntr�;  Rr�;  �r�;  Rr�;  X   JJr�;  G?�      sj^  j  �r�;  h h(h
c__builtin__
__main__
hNN}r�;  Ntr�;  Rr�;  �r�;  Rr�;  (X   ''r�;  G?�-�-�X   NNPr�;  G?���X   INr�;  G?���X   WPr�;  G?��h�hX   VBPr�;  G?��;�;X   WDTr�;  G?��h�hX   CCr�;  G?��h�hhMG?��h�hX   NNr�;  G?���X   CDr�;  G?��h�hX   ``r�;  G?���h�G?���X   VBDr�;  G?��h�hX   POSr�;  G?��h�huX   PRP$r�;  j1
  �r�;  h h(h
c__builtin__
__main__
hNN}r�;  Ntr�;  Rr�;  �r�;  Rr�;  (X   NNSr�;  G?�      X   NNr�;  G?��8�9X   INr�;  G?��q�rX   JJr�;  G?�q�q�X   DTr�;  G?�q�q�h�G?�q�q�uh�j�  �r�;  h h(h
c__builtin__
__main__
hNN}r�;  Ntr�;  Rr�;  �r�;  Rr�;  (X   DTr�;  G?�UUUUUUX   RPr�;  G?�UUUUUUX   INr�;  G?�UUUUUUX   NNPr�;  G?�UUUUUUX   oovr�;  G?�UUUUUUuX   ''r�;  j�  �r�;  h h(h
c__builtin__
__main__
hNN}r�;  Ntr�;  Rr�;  �r�;  Rr�;  (X   INr�;  G?�q�q�h�G?�q�q�X   VBr�;  G?�З�%�	X   WPr�;  G?�����/hX   NNPr�;  G?�����/hX   DTr�;  G?�����/hX   ``r�;  G?�����/huX   ''r�;  j�  �r�;  h h(h
c__builtin__
__main__
hNN}r�;  Ntr�;  Rr�;  �r�;  Rr�;  (X   PRP$r�;  G?��}�pX   ``r�;  G?�tŝ1gX   WPr�;  G?��}�pX   DTr�;  G?�򆼡�(X   VBZr�;  G?�򆼡�(X   NNr <  G?��}�pX   VBPr<  G?��}�pX   RBr<  G?��}�pX   JJr<  G?��}�pX   NNSr<  G?��}�puX   ``r<  j  �r<  h h(h
c__builtin__
__main__
hNN}r<  Ntr<  Rr	<  �r
<  Rr<  (X   RBr<  G?�UUUUUUX   PRPr<  G?�q�q�X   NNPr<  G?�q�q�uX   ``r<  j�  �r<  h h(h
c__builtin__
__main__
hNN}r<  Ntr<  Rr<  �r<  Rr<  (X   DTr<  G?���a|X   VBr<  G?���a{�X   NNSr<  G?���a{�X   PRPr<  G?�{���aX   VBPr<  G?���a{�X   NNr<  G?�{���aX   ''r<  G?���a{�X   NNPr<  G?���a{�X   MDr<  G?���a{�X   VBZr<  G?���a{�h�G?���a{�uX   DTr <  j�  �r!<  h h(h
c__builtin__
__main__
hNN}r"<  Ntr#<  Rr$<  �r%<  Rr&<  (X   VBNr'<  G?�������X   RBr(<  G?�X   INr)<  G?�<<<<<<X   TOr*<  G?�X   PRP$r+<  G?�������X   DTr,<  G?�X   PRPr-<  G?�������hMG?�X   WPr.<  G?�X   NNPr/<  G?�X   VBGr0<  G?�X   NNSr1<  G?�������X   VBDr2<  G?�X   JJr3<  G?�������X   CDr4<  G?�X   WRBr5<  G?�X   NNr6<  G?�uj'<  jL#  �r7<  h h(h
c__builtin__
__main__
hNN}r8<  Ntr9<  Rr:<  �r;<  Rr<<  (X   CDr=<  G?�������X   INr><  G?���Q�X   JJr?<  G?�������X   NNr@<  G?�������X   NNSrA<  G?У�
=p�h�G?�z�G�{X   CCrB<  G?��Q��X   NNPrC<  G?��Q��uX   ``rD<  j�  �rE<  h h(h
c__builtin__
__main__
hNN}rF<  NtrG<  RrH<  �rI<  RrJ<  (X   NNPrK<  G?�      X   ''rL<  G?�UUUUUUX   JJrM<  G?�      X   NNrN<  G?�UUUUUUuX   JJSrO<  j�4  �rP<  h h(h
c__builtin__
__main__
hNN}rQ<  NtrR<  RrS<  �rT<  RrU<  (X   INrV<  G?�t]E�tX   RBrW<  G?�E�t]FX   JJrX<  G?�E�t]FX   NNSrY<  G?�E�t]FX   NNrZ<  G?�E�t]FuX   JJr[<  jf  �r\<  h h(h
c__builtin__
__main__
hNN}r]<  Ntr^<  Rr_<  �r`<  Rra<  (X   NNrb<  G?��q�rX   VBrc<  G?�q�q�X   CDrd<  G?��8�9X   VBPre<  G?�q�q�X   INrf<  G?�q�q�X   DTrg<  G?�UUUUUUX   RBrh<  G?��q�rX   JJri<  G?��q�rX   NNPrj<  G?�q�q�X   VBNrk<  G?�q�q�h�G?�q�q�X   NNSrl<  G?��q�rX   CCrm<  G?�q�q�X   VBZrn<  G?�UUUUUUX   VBGro<  G?�UUUUUUX   ``rp<  G?�UUUUUUuj�  jz8  �rq<  h h(h
c__builtin__
__main__
hNN}rr<  Ntrs<  Rrt<  �ru<  Rrv<  (X   NNPrw<  G?�I$�I$�X   VBNrx<  G?�I$�I$�X   DTry<  G?�UUUUUUX   INrz<  G?�I$�I$�X   NNr{<  G?�a�a�X   JJr|<  G?�UUUUUUX   VBGr}<  G?�I$�I$�h�G?�a�a�X   RBr~<  G?�I$�I$�X   WPr<  G?�a�a�X   PRPr�<  G?�a�a�uX   VBDr�<  j�  �r�<  h h(h
c__builtin__
__main__
hNN}r�<  Ntr�<  Rr�<  �r�<  Rr�<  (X   JJr�<  G?��,��,�X   VBNr�<  G?�AAX   NNr�<  G?�AAX   RBr�<  G?�AAX   NNPSr�<  G?�AAX   NNSr�<  G?�a�a�X   VBr�<  G?�AAX   INr�<  G?�AAX   CDr�<  G?�AAuj�  j�  �r�<  h h(h
c__builtin__
__main__
hNN}r�<  Ntr�<  Rr�<  �r�<  Rr�<  X   VBr�<  G?�      sX   NNSr�<  j�  �r�<  h h(h
c__builtin__
__main__
hNN}r�<  Ntr�<  Rr�<  �r�<  Rr�<  (X   CDr�<  G?�����/hX   PRPr�<  G?�����/hX   JJr�<  G?�q�q�X   INr�<  G?�q�q�X   MDr�<  G?�����/hX   RBr�<  G?�����/hX   VBGr�<  G?�����/hX   VBPr�<  G?�q�q�X   DTr�<  G?�q�q�X   NNPr�<  G?�q�q�h�G?��q�rX   WDTr�<  G?�����/hX   VBZr�<  G?�����/hX   CCr�<  G?�����/hX   JJRr�<  G?�����/huX   PRP$r�<  j�  �r�<  h h(h
c__builtin__
__main__
hNN}r�<  Ntr�<  Rr�<  �r�<  Rr�<  (h�G?�.���/X   INr�<  G?�E�t]Fuj!  j2  �r�<  h h(h
c__builtin__
__main__
hNN}r�<  Ntr�<  Rr�<  �r�<  Rr�<  (X   INr�<  G?�'bv'bvX   RBr�<  G?��;�;X   PRP$r�<  G?��;�;X   DTr�<  G?��;�;X   WRBr�<  G?��;�;h�G?ȝ�؝��X   NNr�<  G?��;�;X   ``r�<  G?��;�;uX   VBNr�<  j+  �r�<  h h(h
c__builtin__
__main__
hNN}r�<  Ntr�<  Rr�<  �r�<  Rr�<  (X   WPr�<  G?�UUUUUUX   VBNr�<  G?�333333X   VBGr�<  G?�X   JJr�<  G?�X   DTr�<  G?�������X   RBr�<  G?�������X   VBZr�<  G?�X   oovr�<  G?�X   INr�<  G?�uX   CCr�<  j�;  �r�<  h h(h
c__builtin__
__main__
hNN}r�<  Ntr�<  Rr�<  �r�<  Rr�<  (X   PRPr�<  G?�X   NNr�<  G?�X   RBr�<  G?�X   JJr�<  G?�������X   INr�<  G?�X   NNPr�<  G?Ɩ�����X   VBNr�<  G?�X   NNSr�<  G?�X   DTr�<  G?�X   JJRr�<  G?�X   VBGr�<  G?�uX   INr�<  j�  �r�<  h h(h
c__builtin__
__main__
hNN}r�<  Ntr�<  Rr�<  �r�<  Rr�<  (X   CDr�<  G?�333333X   VBr�<  G?�333333X   NNPr�<  G?�333333X   WPr�<  G?�������X   RPr�<  G?�333333X   PRPr�<  G?�������X   DTr�<  G?�333333X   INr�<  G?�������X   NNr�<  G?�333333X   RBr�<  G?�      X   JJr�<  G?�      X   VBNr�<  G?�������X   NNSr�<  G?�������uNh2�r�<  h h(h
c__builtin__
__main__
hNN}r�<  Ntr�<  Rr�<  �r�<  Rr�<  (X   INr�<  G?�5�yC^X   NNr�<  G?�1gLY�X   NNSr =  G?�5�yC^X   RBr=  G?�򆼡�(X   TOr=  G?�tŝ1gLX   NNPSr=  G?��}�pX   VBDr=  G?��}�puX   VBPr=  j�  �r=  h h(h
c__builtin__
__main__
hNN}r=  Ntr=  Rr	=  �r
=  Rr=  (X   NNr=  G?��Gq�wX   DTr=  G?��_A}�X   JJRr=  G?��Gq�wX   VBPr=  G?�SYMe5�X   RBr=  G?��_A}�X   JJr=  G?��w�GqX   VBDr=  G?��_A}�X   NNSr=  G?��_A}�X   VBNr=  G?��Gq�wX   VBr=  G?��Gq�wuX   JJSr=  j�  �r=  h h(h
c__builtin__
__main__
hNN}r=  Ntr=  Rr=  �r=  Rr=  (h�G?�      X   NNr=  G?�      X   INr=  G?�      uX   WPr=  ju  �r =  h h(h
c__builtin__
__main__
hNN}r!=  Ntr"=  Rr#=  �r$=  Rr%=  (X   NNr&=  G?ڪ�����h�G?�UUUUUUX   VBGr'=  G?�UUUUUUX   JJr(=  G?�      uX   PRPr)=  j�  �r*=  h h(h
c__builtin__
__main__
hNN}r+=  Ntr,=  Rr-=  �r.=  Rr/=  (X   JJr0=  G?�t]E�tX   NNSr1=  G?�E�t]FX   INr2=  G?�E�t]FX   NNr3=  G?�E�t]Fh�G?�E�t]FuX   NNSr4=  j�  �r5=  h h(h
c__builtin__
__main__
hNN}r6=  Ntr7=  Rr8=  �r9=  Rr:=  (X   NNr;=  G?�;�6w�mX   INr<=  G?�W& �Lh�G?�W& �LAX   CCr==  G?�Ɉ+�WX   RBr>=  G?�Ɉ+�WX   WPr?=  G?�Ɉ+�WX   NNSr@=  G?�W& �LAuX   WPrA=  hM�rB=  h h(h
c__builtin__
__main__
hNN}rC=  NtrD=  RrE=  �rF=  RrG=  (X   INrH=  G?��}�pX   VBGrI=  G?�pG��X   JJrJ=  G?��}�pX   RBrK=  G?�tŝ1gLX   VBDrL=  G?�򆼡�(X   PRPrM=  G?��}�pX   VBZrN=  G?��}�pX   NNrO=  G?��}�pX   WRBrP=  G?��}�puX   WPrQ=  jv  �rR=  h h(h
c__builtin__
__main__
hNN}rS=  NtrT=  RrU=  �rV=  RrW=  (X   RBrX=  G?�I$�I$�h�G?�I$�I$�NG?�m��m��uX   DTrY=  ju  �rZ=  h h(h
c__builtin__
__main__
hNN}r[=  Ntr\=  Rr]=  �r^=  Rr_=  (X   NNr`=  G?�      X   NNPra=  G?�      X   WRBrb=  G?�������X   WPrc=  G?�������X   JJrd=  G?�������X   INre=  G?�������X   DTrf=  G?�������uX   ''rg=  j�2  �rh=  h h(h
c__builtin__
__main__
hNN}ri=  Ntrj=  Rrk=  �rl=  Rrm=  (X   TOrn=  G?�      X   PRP$ro=  G?�      X   PRPrp=  G?�      X   NNSrq=  G?�      NG?�      X   RBrr=  G?�      X   JJrs=  G?�      h�G?�      X   DTrt=  G?�      X   INru=  G?�      uX   NNSrv=  j�  �rw=  h h(h
c__builtin__
__main__
hNN}rx=  Ntry=  Rrz=  �r{=  Rr|=  (X   NNSr}=  G?�      X   JJr~=  G?�      X   NNr=  G?�      X   VBNr�=  G?�      uX   CDr�=  j�4  �r�=  h h(h
c__builtin__
__main__
hNN}r�=  Ntr�=  Rr�=  �r�=  Rr�=  (X   CDr�=  G?��y�zX   WDTr�=  G?�a�a�X   CCr�=  G?�a�a�X   VBZr�=  G?�I$�I$�X   NNPr�=  G?�UUUUUUh�G?�a�a�X   WRBr�=  G?�a�a�X   oovr�=  G?�I$�I$�X   VBNr�=  G?�a�a�X   VBDr�=  G?�a�a�X   JJr�=  G?�a�a�X   RBr�=  G?�a�a�X   NNr�=  G?�a�a�X   DTr�=  G?�a�a�X   ``r�=  G?�a�a�uX   VBZr�=  hM�r�=  h h(h
c__builtin__
__main__
hNN}r�=  Ntr�=  Rr�=  �r�=  Rr�=  (X   WPr�=  G?�I$�I$�X   NNSr�=  G?�A�A�X   WRBr�=  G?��_�_X   PRPr�=  G?�A�A�X   VBNr�=  G?�A�A�X   INr�=  G?�A�A�X   DTr�=  G?�A�A�X   NNPr�=  G?�A�A�X   JJr�=  G?�A�A�X   ``r�=  G?�A�A�uX   PRPr�=  j  �r�=  h h(h
c__builtin__
__main__
hNN}r�=  Ntr�=  Rr�=  �r�=  Rr�=  (X   ''r�=  G?�I$�I$�h�G?�m��m��uj�&  jQ(  �r�=  h h(h
c__builtin__
__main__
hNN}r�=  Ntr�=  Rr�=  �r�=  Rr�=  (X   VBDr�=  G?�UUUUUUX   WDTr�=  G?�      X   NNr�=  G?�UUUUUUh�G?�UUUUUUX   INr�=  G?�UUUUUUX   VBNr�=  G?�UUUUUUX   RBr�=  G?�UUUUUUuX   ''r�=  j�  �r�=  h h(h
c__builtin__
__main__
hNN}r�=  Ntr�=  Rr�=  �r�=  Rr�=  (X   NNPr�=  G?�UUUUUUX   VBZr�=  G?�UUUUUUX   VBDr�=  G?ʪ�����X   MDr�=  G?�UUUUUUX   VBPr�=  G?�UUUUUUuX   WRBr�=  j�  �r�=  h h(h
c__builtin__
__main__
hNN}r�=  Ntr�=  Rr�=  �r�=  Rr�=  (X   VBDr�=  G?�      X   VBZr�=  G?�      X   NNr�=  G?�      X   MDr�=  G?�      uX   DTr�=  j�  �r�=  h h(h
c__builtin__
__main__
hNN}r�=  Ntr�=  Rr�=  �r�=  Rr�=  (X   VBr�=  G?�����/hX   INr�=  G?�����/hh�G?�q�q�uX   CDr�=  j5  �r�=  h h(h
c__builtin__
__main__
hNN}r�=  Ntr�=  Rr�=  �r�=  Rr�=  (X   VBr�=  G?�E�t]X   RBr�=  G?�E�t]FuX   VBDr�=  hM�r�=  h h(h
c__builtin__
__main__
hNN}r�=  Ntr�=  Rr�=  �r�=  Rr�=  (X   WRBr�=  G?�q�q�X   JJr�=  G?���<�XX   WPr�=  G?��<�X~X   ``r�=  G?���<�XX   DTr�=  G?�����/hX   VBDr�=  G?�����/hX   CCr�=  G?���<�XX   INr�=  G?�����/hX   VBGr�=  G?�H�����X   NNPr�=  G?�����/hX   CDr�=  G?�H�����X   NNr�=  G?�����/hX   WDTr�=  G?�H�����X   RBr�=  G?�H�����X   TOr�=  G?�H�����X   VBr�=  G?�H�����X   PRPr�=  G?�����/huX   JJr�=  j�  �r�=  h h(h
c__builtin__
__main__
hNN}r�=  Ntr�=  Rr >  �r>  Rr>  (X   VBZr>  G?��m��m�X   VBDr>  G?�I$�I$�X   NNr>  G?�I$�I$�X   MDr>  G?�I$�I$�X   VBPr>  G?�I$�I$�uX   NNPSr>  j3  �r	>  h h(h
c__builtin__
__main__
hNN}r
>  Ntr>  Rr>  �r>  Rr>  (X   INr>  G?�      X   MDr>  G?�������X   NNPr>  G?ə�����X   VBPr>  G?�������h�G?�      X   VBDr>  G?�������uX   CDr>  j�  �r>  h h(h
c__builtin__
__main__
hNN}r>  Ntr>  Rr>  �r>  Rr>  (X   NNr>  G?��a���X   VBDr>  G?��A)��X   INr>  G?��a���X   VBNr>  G?��a���X   CDr>  G?��A)��X   JJr >  G?�Jy��JX   VBZr!>  G?��a���X   RBr">  G?��A)��h�G?�E�t]FX   VBr#>  G?��a���X   WRBr$>  G?��A)��X   VBPr%>  G?�E�t]FX   VBGr&>  G?��A)��X   NNSr'>  G?��A)��uX   ''r(>  j/  �r)>  h h(h
c__builtin__
__main__
hNN}r*>  Ntr+>  Rr,>  �r->  Rr.>  (X   VBr/>  G?�'bv'bvX   RBr0>  G?ñ;�;X   DTr1>  G?ñ;�;uj�"  j�"  �r2>  h h(h
c__builtin__
__main__
hNN}r3>  Ntr4>  Rr5>  �r6>  Rr7>  (X   JJr8>  G?�UUUUUUX   NNSr9>  G?�X   NNr:>  G?�X   JJSr;>  G?�uX   VBr<>  j2  �r=>  h h(h
c__builtin__
__main__
hNN}r>>  Ntr?>  Rr@>  �rA>  RrB>  (X   WPrC>  G?�I$�I$�X   JJrD>  G?�m��m��X   VBNrE>  G?�m��m��X   INrF>  G?�m��m��X   DTrG>  G?�m��m��X   PRP$rH>  G?�I$�I$�X   NNSrI>  G?�m��m��X   TOrJ>  G?�I$�I$�X   PRPrK>  G?�I$�I$�X   NNPSrL>  G?�I$�I$�uhMj�"  �rM>  h h(h
c__builtin__
__main__
hNN}rN>  NtrO>  RrP>  �rQ>  RrR>  (X   WRBrS>  G?��!B�X   CDrT>  G?��!B�X   VBNrU>  G?��1�c�X   NNSrV>  G?��9�s��X   WPrW>  G?��!B�X   PRPrX>  G?��1�c�X   PRP$rY>  G?��1�c�X   NNrZ>  G?��)JR��X   INr[>  G?ĥ)JR��X   JJr\>  G?��1�c�X   JJSr]>  G?��!B�X   DTr^>  G?��1�c�X   oovr_>  G?��!B�X   WDTr`>  G?��!B�X   NNPra>  G?��!B�X   TOrb>  G?��1�c�X   RBrc>  G?��!B�uNh3�rd>  h h(h
c__builtin__
__main__
hNN}re>  Ntrf>  Rrg>  �rh>  Rri>  (X   JJRrj>  G?�a�AvX   DTrk>  G?�UUUUUUX   NNSrl>  G?���z�^�X   PRPrm>  G?����X   JJrn>  G?�������X   VBDro>  G?���+@X   NNrp>  G?�a�AvX   NNPrq>  G?����X   WPrr>  G?���+@X   VBGrs>  G?���+@X   CDrt>  G?����X   PRP$ru>  G?���+@X   NNPSrv>  G?���+@X   JJSrw>  G?���+@uX   oovrx>  j�  �ry>  h h(h
c__builtin__
__main__
hNN}rz>  Ntr{>  Rr|>  �r}>  Rr~>  (X   JJr>  G?�I$�I$�X   DTr�>  G?��m��m�X   TOr�>  G?�I$�I$�X   PRP$r�>  G?�m��m��X   oovr�>  G?�I$�I$�h�G?�m��m��X   INr�>  G?�I$�I$�X   VBNr�>  G?�I$�I$�X   NNSr�>  G?�I$�I$�X   NNr�>  G?�I$�I$�uX   JJSr�>  j  �r�>  h h(h
c__builtin__
__main__
hNN}r�>  Ntr�>  Rr�>  �r�>  Rr�>  (X   CCr�>  G?�      X   NNPr�>  G?�      X   DTr�>  G?�      X   INr�>  G?�      uX   ``r�>  j  �r�>  h h(h
c__builtin__
__main__
hNN}r�>  Ntr�>  Rr�>  �r�>  Rr�>  (X   ''r�>  G?��i�XGX   VBNr�>  G?�{���aX   INr�>  G?�{���aX   JJr�>  G?���a{�h�G?�{���aX   NNr�>  G?���a{�uj�>  j�6  �r�>  h h(h
c__builtin__
__main__
hNN}r�>  Ntr�>  Rr�>  �r�>  Rr�>  (X   VBPr�>  G?�q�q�h�G?�EQEQX   INr�>  G?�AAX   TOr�>  G?�QEQEX   MDr�>  G?�AAX   VBDr�>  G?�QEQEX   NNr�>  G?�AAX   VBNr�>  G?�AAX   JJr�>  G?�AAX   VBGr�>  G?�AAX   VBr�>  G?�AAX   RBr�>  G?�AAujT  jD:  �r�>  h h(h
c__builtin__
__main__
hNN}r�>  Ntr�>  Rr�>  �r�>  Rr�>  (X   NNr�>  G?�      X   NNSr�>  G?��8�9h�G?��8�9X   VBr�>  G?�q�q�X   VBGr�>  G?�q�q�X   oovr�>  G?�q�q�X   NNPr�>  G?�UUUUUUX   TOr�>  G?�q�q�X   NNPSr�>  G?�q�q�uX   VBNr�>  j�  �r�>  h h(h
c__builtin__
__main__
hNN}r�>  Ntr�>  Rr�>  �r�>  Rr�>  (X   RBr�>  G?�i��i��X   NNr�>  G?�AAX   JJr�>  G?�AAX   TOr�>  G?�a�a�X   WRBr�>  G?�AAX   INr�>  G?�q�q�X   CDr�>  G?�a�a�h�G?�AAX   DTr�>  G?�AAhMG?�AAX   VBPr�>  G?�AAX   oovr�>  G?�AAX   PRPr�>  G?�AAX   ``r�>  G?�a�a�uj�%  hM�r�>  h h(h
c__builtin__
__main__
hNN}r�>  Ntr�>  Rr�>  �r�>  Rr�>  (X   NNSr�>  G?�X   PRPr�>  G?�������X   VBGr�>  G?�������X   WPr�>  G?�X   VBPr�>  G?�X   RBr�>  G?�������X   VBNr�>  G?�X   WRBr�>  G?�X   CCr�>  G?�������X   NNPr�>  G?�X   INr�>  G?�X   NNr�>  G?�uX   CDr�>  j�
  �r�>  h h(h
c__builtin__
__main__
hNN}r�>  Ntr�>  Rr�>  �r�>  Rr�>  (h�G?̨�1��X   NNr�>  G?�&5~��X   JJr�>  G?���@�X   NNPr�>  G?��vr�zX   CDr�>  G?��1��gX   JJSr�>  G?���@�X   NNSr�>  G?��1��gX   RBSr�>  G?���@�X   INr�>  G?��1��guhMj�"  �r�>  h h(h
c__builtin__
__main__
hNN}r�>  Ntr�>  Rr�>  �r�>  Rr�>  (X   VBPr�>  G?�gȦ�}X   VBZr�>  G?��>E0oX   MDr�>  G?�7Y�)�vX   VBDr�>  G?�"�7Y�*X   RBr�>  G?���ϑLuX   JJRr�>  jG/  �r�>  h h(h
c__builtin__
__main__
hNN}r�>  Ntr ?  Rr?  �r?  Rr?  (X   DTr?  G?�I$�I%X   NNPr?  G?�m��m��X   oovr?  G?�I$�I$�uX   JJRr?  jN1  �r?  h h(h
c__builtin__
__main__
hNN}r	?  Ntr
?  Rr?  �r?  Rr?  (X   INr?  G?�      X   DTr?  G?�      uX   CDr?  j�
  �r?  h h(h
c__builtin__
__main__
hNN}r?  Ntr?  Rr?  �r?  Rr?  (X   NNPr?  G?�R�+x�X   CDr?  G?��+x�5"X   NNSr?  G?�&�9�V�X   TOr?  G?�R�+x�X   NNr?  G?��+x�5"X   INr?  G?��+x�5"X   WPr?  G?�R�+x�X   DTr?  G?ż`����X   PRP$r?  G?�R�+x�X   VBGr ?  G?�R�+x�h�G?�R�+x�uX   NNPSr!?  j  �r"?  h h(h
c__builtin__
__main__
hNN}r#?  Ntr$?  Rr%?  �r&?  Rr'?  (X   NNPr(?  G?�q�q�h�G?�UUUUUUX   NNSr)?  G?�q�q�X   JJr*?  G?�q�q�uX   CCr+?  j�  �r,?  h h(h
c__builtin__
__main__
hNN}r-?  Ntr.?  Rr/?  �r0?  Rr1?  (h�G?�I$�I$�X   VBr2?  G?��m��m�X   WDTr3?  G?�I$�I$�X   WPr4?  G?�I$�I$�X   DTr5?  G?�m��m��uX   RPr6?  j  �r7?  h h(h
c__builtin__
__main__
hNN}r8?  Ntr9?  Rr:?  �r;?  Rr<?  (X   VBr=?  G?�      X   RBr>?  G?�UUUUUUX   VBDr??  G?�UUUUUUX   VBGr@?  G?�UUUUUUuX   VBPrA?  j
  �rB?  h h(h
c__builtin__
__main__
hNN}rC?  NtrD?  RrE?  �rF?  RrG?  (X   RBrH?  G?�      X   DTrI?  G?�������X   VBrJ?  G?ᙙ����X   RBSrK?  G?�������uX   VBGrL?  jG  �rM?  h h(h
c__builtin__
__main__
hNN}rN?  NtrO?  RrP?  �rQ?  RrR?  (X   VBrS?  G?↼��(lX   RBrT?  G?�5�yC^X   DTrU?  G?�5�yC^X   PRPrV?  G?�򆼡�(uX   INrW?  j�  �rX?  h h(h
c__builtin__
__main__
hNN}rY?  NtrZ?  Rr[?  �r\?  Rr]?  (X   VBr^?  G?��q�rh�G?�q�q�hMG?�q�q�X   RBr_?  G?�q�q�X   PRPr`?  G?�q�q�uX   VBGra?  j�&  �rb?  h h(h
c__builtin__
__main__
hNN}rc?  Ntrd?  Rre?  �rf?  Rrg?  (X   NNSrh?  G?�B�Y!dX   INri?  G?вB�YX   NNrj?  G?��B�YX   JJrk?  G?��zoM�X   VBNrl?  G?��B�Yh�G?�B�Y!dX   CCrm?  G?�B�Y!dX   NNPSrn?  G?�B�Y!dhMG?�B�Y!dX   TOro?  G?�B�Y!dX   DTrp?  G?�B�Y!duX   WDTrq?  j4  �rr?  h h(h
c__builtin__
__main__
hNN}rs?  Ntrt?  Rru?  �rv?  Rrw?  (X   NNSrx?  G?�q�q�X   NNry?  G?�UUUUUUX   VBPrz?  G?�q�q�X   VBDr{?  G?�q�q�uX   JJr|?  j  �r}?  h h(h
c__builtin__
__main__
hNN}r~?  Ntr?  Rr�?  �r�?  Rr�?  (h�G?З�%�	{X   NNr�?  G?״%�	{BX   NNSr�?  G?�����/hX   DTr�?  G?�����/hX   JJSr�?  G?�����/hX   JJr�?  G?�����/huX   VBZr�?  j�  �r�?  h h(h
c__builtin__
__main__
hNN}r�?  Ntr�?  Rr�?  �r�?  Rr�?  (X   NNPr�?  G?ə�����h�G?�X   oovr�?  G?�X   VBr�?  G?�X   VBGr�?  G?�X   NNr�?  G?�uh�j�  �r�?  h h(h
c__builtin__
__main__
hNN}r�?  Ntr�?  Rr�?  �r�?  Rr�?  (X   NNPr�?  G?ñ;�;X   NNr�?  G?ñ;�;X   JJr�?  G?ñ;�;X   DTr�?  G?ñ;�;NG?؝�؝��uh�j�  �r�?  h h(h
c__builtin__
__main__
hNN}r�?  Ntr�?  Rr�?  �r�?  Rr�?  (X   DTr�?  G?�      X   CDr�?  G?�������X   NNPr�?  G?�      X   JJr�?  G?�������h�G?�������X   NNr�?  G?�������X   RBr�?  G?�������uX   VBDr�?  j�  �r�?  h h(h
c__builtin__
__main__
hNN}r�?  Ntr�?  Rr�?  �r�?  Rr�?  (X   PRP$r�?  G?�UUUUUUX   DTr�?  G?�      X   RBr�?  G?�UUUUUUX   JJr�?  G?�      X   INr�?  G?�UUUUUUuX   TOr�?  j�*  �r�?  h h(h
c__builtin__
__main__
hNN}r�?  Ntr�?  Rr�?  �r�?  Rr�?  (X   VBGr�?  G?ñ;�;X   INr�?  G?�;�;�X   RBr�?  G?ñ;�;X   VBr�?  G?ñ;�;uX   JJSr�?  j  �r�?  h h(h
c__builtin__
__main__
hNN}r�?  Ntr�?  Rr�?  �r�?  Rr�?  (X   RBSr�?  G?�m��m��X   JJSr�?  G?�m��m��X   VBr�?  G?�I$�I$�X   JJr�?  G?�m��m��X   RBr�?  G?�m��m��uj  j�?  �r�?  h h(h
c__builtin__
__main__
hNN}r�?  Ntr�?  Rr�?  �r�?  Rr�?  (X   JJr�?  G?陙����X   RBr�?  G?ə�����uX   CCr�?  j�?  �r�?  h h(h
c__builtin__
__main__
hNN}r�?  Ntr�?  Rr�?  �r�?  Rr�?  (X   NNSr�?  G?��8�9X   NNr�?  G?�UUUUUUX   INr�?  G?�UUUUUUh�G?�q�q�X   TOr�?  G?�q�q�X   JJr�?  G?�q�q�hMG?�q�q�X   ''r�?  G?�q�q�uX   CCr�?  j�1  �r�?  h h(h
c__builtin__
__main__
hNN}r�?  Ntr�?  Rr�?  �r�?  Rr�?  (X   INr�?  G?����� h�G?ũZ��Z�X   NNPr�?  G?��;�;X   VBDr�?  G?����� hMG?��;�;X   VBPr�?  G?����� X   VBNr�?  G?��z�zX   MDr�?  G?����� X   NNSr�?  G?��z�zX   VBGr�?  G?����� X   NNPSr�?  G?����� X   VBr�?  G?����� X   CCr�?  G?����� X   RBr�?  G?����� X   TOr�?  G?����� uX   WDTr�?  j!:  �r�?  h h(h
c__builtin__
__main__
hNN}r�?  Ntr�?  Rr�?  �r�?  Rr�?  (X   PRP$r�?  G?�UUUUUUX   NNr�?  G?�UUUUUUuX   PRPr�?  jH$  �r @  h h(h
c__builtin__
__main__
hNN}r@  Ntr@  Rr@  �r@  Rr@  (X   NNSr@  G?�X   JJr@  G?�X   PRPr@  G?�ZZZZZZX   NNr	@  G?�X   DTr
@  G?�X   TOr@  G?�uX   WDTr@  j�  �r@  h h(h
c__builtin__
__main__
hNN}r@  Ntr@  Rr@  �r@  Rr@  (X   NNr@  G?�m��m��X   VBZr@  G?�I$�I$�X   JJr@  G?�I$�I$�ujk  j�8  �r@  h h(h
c__builtin__
__main__
hNN}r@  Ntr@  Rr@  �r@  Rr@  (X   VBPr@  G?��SYMe6h�G?�YMe5��X   VBr@  G?��_A}�X   NNr@  G?��_A}�X   CCr@  G?��_A}�X   MDr @  G?��_A}�X   VBGr!@  G?��_A}�X   VBDr"@  G?��Gq�wX   INr#@  G?��w�GquX   ''r$@  j�  �r%@  h h(h
c__builtin__
__main__
hNN}r&@  Ntr'@  Rr(@  �r)@  Rr*@  (X   VBNr+@  G?�X   TOr,@  G?ٙ�����X   NNr-@  G?ə�����X   INr.@  G?�X   RBr/@  G?�uX   VBNr0@  j�  �r1@  h h(h
c__builtin__
__main__
hNN}r2@  Ntr3@  Rr4@  �r5@  Rr6@  (X   DTr7@  G?�UUUUUUX   NNPr8@  G?�UUUUUUh�G?�UUUUUUX   NNr9@  G?�      X   VBr:@  G?�UUUUUUX   NNSr;@  G?�UUUUUUX   JJr<@  G?�      X   oovr=@  G?�UUUUUUX   VBPr>@  G?�UUUUUUuNh4�r?@  h h(h
c__builtin__
__main__
hNN}r@@  NtrA@  RrB@  �rC@  RrD@  (X   PRPrE@  G?�4[_uX   DTrF@  G?�<��N	X   VBGrG@  G?�[_u'X   NNrH@  G?�[_u'X   NNSrI@  G?��I�A�X   CDrJ@  G?���/��X   VBrK@  G?�[_u'X   JJrL@  G?�_u'WX   NNPrM@  G?����Rp�X   MDrN@  G?�[_u'X   RBrO@  G?���/��uX   JJRrP@  j2  �rQ@  h h(h
c__builtin__
__main__
hNN}rR@  NtrS@  RrT@  �rU@  RrV@  (X   NNrW@  G?��;�;X   JJRrX@  G?�؝�؞X   JJrY@  G?��;�;X   oovrZ@  G?ȝ�؝��X   NNPr[@  G?��؝�؞uX   WRBr\@  j/   �r]@  h h(h
c__builtin__
__main__
hNN}r^@  Ntr_@  Rr`@  �ra@  Rrb@  (X   WRBrc@  G?�'bv'bvX   WPrd@  G?ñ;�;X   INre@  G?ñ;�;uj/   jc@  �rf@  h h(h
c__builtin__
__main__
hNN}rg@  Ntrh@  Rri@  �rj@  Rrk@  (X   PRPrl@  G?�q�q�X   JJrm@  G?�UUUUUUh�G?�����/hX   RBrn@  G?�q�q�X   DTro@  G?�����/hX   VBDrp@  G?�����/X   CCrq@  G?�����/hX   VBZrr@  G?�q�q�NG?�����/hX   VBPrs@  G?�����/hX   NNrt@  G?�����/hX   MDru@  G?�q�q�uX   VBGrv@  jH  �rw@  h h(h
c__builtin__
__main__
hNN}rx@  Ntry@  Rrz@  �r{@  Rr|@  (X   VBNr}@  G?��1�c�X   INr~@  G?��1�c�h�G?��!B�X   JJRr@  G?��!B�X   TOr�@  G?��1�c�X   DTr�@  G?��!B�X   NNPr�@  G?��1�c�X   WPr�@  G?��1�c�X   NNSr�@  G?ĥ)JR��uX   ''r�@  j3  �r�@  h h(h
c__builtin__
__main__
hNN}r�@  Ntr�@  Rr�@  �r�@  Rr�@  (X   NNr�@  G?䴴����X   JJr�@  G?�X   NNPr�@  G?�uhMj9  �r�@  h h(h
c__builtin__
__main__
hNN}r�@  Ntr�@  Rr�@  �r�@  Rr�@  (X   NNr�@  G?�UUUUUUX   VBPr�@  G?�      X   VBDr�@  G?�      X   MDr�@  G?�UUUUUUhMG?�      X   CDr�@  G?�      h�G?ª�����X   NNSr�@  G?�UUUUUUX   VBZr�@  G?�      X   JJr�@  G?�UUUUUUX   CCr�@  G?�UUUUUUX   NNPr�@  G?�UUUUUUuhMj�  �r�@  h h(h
c__builtin__
__main__
hNN}r�@  Ntr�@  Rr�@  �r�@  Rr�@  (X   VBGr�@  G?������X   VBr�@  G?ډ]��ډX   RBr�@  G?��Q+��X   DTr�@  G?�81�8X   PRP$r�@  G?������X   PRPr�@  G?�ډ]���X   NNSr�@  G?��Q+��X   MDr�@  G?������uj�  j�@  �r�@  h h(h
c__builtin__
__main__
hNN}r�@  Ntr�@  Rr�@  �r�@  Rr�@  (X   INr�@  G?�I$�I$�X   NNPr�@  G?�m��m��X   NNSr�@  G?�m��m��X   RBr�@  G?�I$�I$�X   VBr�@  G?�I$�I$�X   TOr�@  G?�I$�I$�X   DTr�@  G?�m��m��X   NNr�@  G?�I$�I$�X   JJr�@  G?�I$�I$�uX   WDTr�@  ji*  �r�@  h h(h
c__builtin__
__main__
hNN}r�@  Ntr�@  Rr�@  �r�@  Rr�@  (X   VBDr�@  G?�UUUUUUX   DTr�@  G?�UUUUUUX   VBr�@  G?�UUUUUUuji*  j�@  �r�@  h h(h
c__builtin__
__main__
hNN}r�@  Ntr�@  Rr�@  �r�@  Rr�@  (X   VBNr�@  G?�      X   NNSr�@  G?�      uX   NNSr�@  N�r�@  h h(h
c__builtin__
__main__
hNN}r�@  Ntr�@  Rr�@  �r�@  Rr�@  NG?�      sX   MDr�@  hM�r�@  h h(h
c__builtin__
__main__
hNN}r�@  Ntr�@  Rr�@  �r�@  Rr�@  (X   INr�@  G?�UUUUUUX   CCr�@  G?�UUUUUUX   VBr�@  G?�UUUUUUuX   POSr�@  j�0  �r�@  h h(h
c__builtin__
__main__
hNN}r�@  Ntr�@  Rr�@  �r�@  Rr�@  (X   INr�@  G?�{���aX   RBr�@  G?�{���aX   oovr�@  G?���a{�X   RPr�@  G?���a{�X   WPr�@  G?���a{�X   DTr�@  G?���a|X   VBNr�@  G?ѧ�a{�X   NNr�@  G?���a{�X   JJr�@  G?���a{�uX   PRP$r�@  j�  �r�@  h h(h
c__builtin__
__main__
hNN}r�@  Ntr�@  Rr�@  �r�@  Rr�@  (X   NNPr�@  G?�      X   PRP$r�@  G?�      uj�  j�%  �r�@  h h(h
c__builtin__
__main__
hNN}r�@  Ntr�@  Rr�@  �r�@  Rr�@  (X   POSr�@  G?��B�YX   RBr�@  G?�B�Y!dh�G?�B�Y!dX   CCr A  G?�B�Y!dX   NNPrA  G?вB�YX   NNSrA  G?�B�Y!dX   NNrA  G?�B�Y!duX   VBNrA  j_  �rA  h h(h
c__builtin__
__main__
hNN}rA  NtrA  RrA  �r	A  Rr
A  (X   INrA  G?�UUUUUUX   VBDrA  G?�q�q�X   CCrA  G?�q�q�X   oovrA  G?�q�q�uX   ``rA  j�  �rA  h h(h
c__builtin__
__main__
hNN}rA  NtrA  RrA  �rA  RrA  X   NNrA  G?�      sh�j�  �rA  h h(h
c__builtin__
__main__
hNN}rA  NtrA  RrA  �rA  RrA  h�G?�      sX   NNPSrA  j3  �rA  h h(h
c__builtin__
__main__
hNN}rA  Ntr A  Rr!A  �r"A  Rr#A  (X   VBDr$A  G?�      X   NNr%A  G?�      uX   NNPSr&A  j3  �r'A  h h(h
c__builtin__
__main__
hNN}r(A  Ntr)A  Rr*A  �r+A  Rr,A  X   INr-A  G?�      sj6  j�8  �r.A  h h(h
c__builtin__
__main__
hNN}r/A  Ntr0A  Rr1A  �r2A  Rr3A  (X   VBPr4A  G?ĥ)JR��X   VBDr5A  G?�c�1�h�G?��!B�X   RBr6A  G?��!B�X   NNr7A  G?��!B�X   VBZr8A  G?��1�c�uX   VBr9A  j5  �r:A  h h(h
c__builtin__
__main__
hNN}r;A  Ntr<A  Rr=A  �r>A  Rr?A  (X   JJr@A  G?�      X   CCrAA  G?�UUUUUUX   NNSrBA  G?�      X   RBrCA  G?�      X   ``rDA  G?�UUUUUUX   DTrEA  G?�UUUUUUX   oovrFA  G?�UUUUUUX   NNPrGA  G?�UUUUUUX   CDrHA  G?�UUUUUUX   ''rIA  G?�UUUUUUX   INrJA  G?�      X   NNrKA  G?�UUUUUUhMG?�UUUUUUh�G?�      X   VBGrLA  G?�UUUUUUX   VBPrMA  G?�      X   VBDrNA  G?�UUUUUUuhMj�"  �rOA  h h(h
c__builtin__
__main__
hNN}rPA  NtrQA  RrRA  �rSA  RrTA  (X   DTrUA  G?�������X   CCrVA  G?�333333X   VBDrWA  G?�333333hMG?�      X   INrXA  G?�������X   WPrYA  G?�������uj�"  jUA  �rZA  h h(h
c__builtin__
__main__
hNN}r[A  Ntr\A  Rr]A  �r^A  Rr_A  (X   VBPr`A  G?�UUUUUUX   NNraA  G?�UUUUUUX   VBDrbA  G?�UUUUUUX   VBGrcA  G?�UUUUUUX   NNPrdA  G?�      X   JJreA  G?ʪ�����X   INrfA  G?�UUUUUUuj�  jR  �rgA  h h(h
c__builtin__
__main__
hNN}rhA  NtriA  RrjA  �rkA  RrlA  (X   oovrmA  G?�E�t]FX   VBrnA  G?�E�t]FX   NNProA  G?�E�t]Fh�G?�t]E�tuX   POSrpA  jU5  �rqA  h h(h
c__builtin__
__main__
hNN}rrA  NtrsA  RrtA  �ruA  RrvA  (X   VBrwA  G?��m��m�X   DTrxA  G?�I$�I$�X   WRBryA  G?�I$�I$�uX   MDrzA  j�  �r{A  h h(h
c__builtin__
__main__
hNN}r|A  Ntr}A  Rr~A  �rA  Rr�A  (X   JJr�A  G?�UUUUUUX   VBNr�A  G?�      h�G?�      X   VBr�A  G?�UUUUUUX   NNSr�A  G?�UUUUUUuX   RBSr�A  j]  �r�A  h h(h
c__builtin__
__main__
hNN}r�A  Ntr�A  Rr�A  �r�A  Rr�A  (X   DTr�A  G?�UUUUUUX   VBr�A  G?�UUUUUUX   VBGr�A  G?�UUUUUUuX   ''r�A  j�  �r�A  h h(h
c__builtin__
__main__
hNN}r�A  Ntr�A  Rr�A  �r�A  Rr�A  (X   CCr�A  G?�      h�G?�      uh�j3  �r�A  h h(h
c__builtin__
__main__
hNN}r�A  Ntr�A  Rr�A  �r�A  Rr�A  (X   TOr�A  G?ə�����X   NNr�A  G?�X   DTr�A  G?ə�����X   NNPr�A  G?�X   PRPr�A  G?ə�����X   INr�A  G?�uX   POSr�A  j�  �r�A  h h(h
c__builtin__
__main__
hNN}r�A  Ntr�A  Rr�A  �r�A  Rr�A  (X   NNr�A  G?�333333h�G?ə�����X   RBr�A  G?�333333X   VBNr�A  G?ə�����uX   NNPSr�A  j3  �r�A  h h(h
c__builtin__
__main__
hNN}r�A  Ntr�A  Rr�A  �r�A  Rr�A  (X   INr�A  G?�������X   NNr�A  G?�h�G?�X   VBr�A  G?�X   PRPr�A  G?�X   NNSr�A  G?�X   NNPSr�A  G?�X   VBZr�A  G?�X   NNPr�A  G?�X   TOr�A  G?�X   CCr�A  G?�X   JJr�A  G?�uX   INr�A  jC  �r�A  h h(h
c__builtin__
__main__
hNN}r�A  Ntr�A  Rr�A  �r�A  Rr�A  (X   NNSr�A  G?��_A}�X   NNPr�A  G?��w�GqX   INr�A  G?��SYMe6X   VBGr�A  G?��Gq�wX   NNr�A  G?��Gq�wX   RBr�A  G?��_A}�X   JJr�A  G?��k)���X   PRPr�A  G?��Gq�wX   PRP$r�A  G?��Gq�wX   RPr�A  G?��_A}�X   WRBr�A  G?��_A}�X   DTr�A  G?��SYMe6X   WPr�A  G?��_A}�X   VBDr�A  G?��_A}�X   CDr�A  G?��_A}�X   VBr�A  G?��_A}�X   VBNr�A  G?��w�GqX   WDTr�A  G?��_A}�X   JJRr�A  G?��_A}�h�G?��_A}�X   ``r�A  G?��_A}�uX   VBPr�A  j   �r�A  h h(h
c__builtin__
__main__
hNN}r�A  Ntr�A  Rr�A  �r�A  Rr�A  (X   DTr�A  G?��l�lX   NNSr�A  G?�X   NNPr�A  G?�q�q�X   RBr�A  G?�X   JJr�A  G?�UUUUUUX   VBr�A  G?��l�lX   NNr�A  G?�X   TOr�A  G?��l�lh�G?��l�lX   JJRr�A  G?��l�luj/  jG
  �r�A  h h(h
c__builtin__
__main__
hNN}r�A  Ntr�A  Rr�A  �r�A  Rr�A  (X   JJr�A  G?�m��m��X   NNr�A  G?�I$�I$�h�G?�I$�I$�X   TOr�A  G?�I$�I$�X   RBr�A  G?�I$�I$�X   DTr�A  G?�m��m��uX   JJRr�A  jH/  �r�A  h h(h
c__builtin__
__main__
hNN}r�A  Ntr�A  Rr�A  �r�A  Rr�A  (X   DTr�A  G?�UUUUUUX   NNPr�A  G?�UUUUUUX   NNSr�A  G?�UUUUUUuX   CCr�A  jE&  �r B  h h(h
c__builtin__
__main__
hNN}rB  NtrB  RrB  �rB  RrB  (X   RBrB  G?��!B�X   ``rB  G?��!B�X   JJrB  G?��!B�X   DTr	B  G?��9�s��X   INr
B  G?��1�c�X   PRPrB  G?��)JR��X   oovrB  G?��!B�X   VBrB  G?��!B�X   NNrB  G?��)JR��X   VBNrB  G?��)JR��X   TOrB  G?��1�c�X   NNSrB  G?��!B�X   PRP$rB  G?��!B�uX   VBDrB  j�  �rB  h h(h
c__builtin__
__main__
hNN}rB  NtrB  RrB  �rB  RrB  (X   VBrB  G?�      X   RBrB  G?�UUUUUUX   DTrB  G?�      X   TOrB  G?�UUUUUUX   JJrB  G?�UUUUUUX   CDrB  G?�      uX   WRBr B  jR  �r!B  h h(h
c__builtin__
__main__
hNN}r"B  Ntr#B  Rr$B  �r%B  Rr&B  (X   VBZr'B  G?�UUUUUUX   VBPr(B  G?״%�	{BX   NNSr)B  G?�����/hX   DTr*B  G?�����/hX   VBDr+B  G?�����/hX   INr,B  G?�����/huX   oovr-B  j�5  �r.B  h h(h
c__builtin__
__main__
hNN}r/B  Ntr0B  Rr1B  �r2B  Rr3B  (h�G?ñ;�;X   VBZr4B  G?��;�;uX   VBDr5B  j�  �r6B  h h(h
c__builtin__
__main__
hNN}r7B  Ntr8B  Rr9B  �r:B  Rr;B  (X   NNr<B  G?��t]E�h�G?�E�t]FX   VBr=B  G?�      X   JJr>B  G?�E�t]FX   CCr?B  G?�E�t]FX   TOr@B  G?�t]E�tX   VBGrAB  G?�E�t]X   RBrBB  G?�E�t]FX   VBNrCB  G?�t]E�tX   DTrDB  G?�t]E�tX   NNSrEB  G?�E�t]FX   ''rFB  G?�E�t]FX   INrGB  G?�E�t]FuX   NNPSrHB  N�rIB  h h(h
c__builtin__
__main__
hNN}rJB  NtrKB  RrLB  �rMB  RrNB  NG?�      sX   VBGrOB  j�  �rPB  h h(h
c__builtin__
__main__
hNN}rQB  NtrRB  RrSB  �rTB  RrUB  (X   JJrVB  G?�������X   INrWB  G?�������X   NNrXB  G?�������X   POSrYB  G?�������X   CCrZB  G?�������X   RBr[B  G?�333333X   NNSr\B  G?�������X   VBNr]B  G?�333333X   DTr^B  G?�������X   ``r_B  G?�������X   PRP$r`B  G?�333333uj�  hM�raB  h h(h
c__builtin__
__main__
hNN}rbB  NtrcB  RrdB  �reB  RrfB  (X   NNPrgB  G?�������X   INrhB  G?�X   WPriB  G?ə�����X   WRBrjB  G?�������X   VBDrkB  G?�X   CCrlB  G?�������X   JJrmB  G?�������X   DTrnB  G?�������X   WDTroB  G?�������uX   JJRrpB  jG2  �rqB  h h(h
c__builtin__
__main__
hNN}rrB  NtrsB  RrtB  �ruB  RrvB  (X   NNPrwB  G?�UUUUUUX   INrxB  G?�      X   VBNryB  G?�UUUUUUuX   NNrzB  j  �r{B  h h(h
c__builtin__
__main__
hNN}r|B  Ntr}B  Rr~B  �rB  Rr�B  (h�G?�UUUUUUhMG?�UUUUUUX   TOr�B  G?�      X   MDr�B  G?�      X   VBPr�B  G?�      X   INr�B  G?�UUUUUUX   VBDr�B  G?�UUUUUUX   JJr�B  G?�UUUUUUuX   POSr�B  j�  �r�B  h h(h
c__builtin__
__main__
hNN}r�B  Ntr�B  Rr�B  �r�B  Rr�B  (X   DTr�B  G?�333333X   VBNr�B  G?ٙ�����X   VBr�B  G?�������X   NNPr�B  G?�������X   RBr�B  G?�������uX   DTr�B  j!  �r�B  h h(h
c__builtin__
__main__
hNN}r�B  Ntr�B  Rr�B  �r�B  Rr�B  (X   POSr�B  G?�I$�I$�X   NNr�B  G?��m��m�uX   INr�B  j�  �r�B  h h(h
c__builtin__
__main__
hNN}r�B  Ntr�B  Rr�B  �r�B  Rr�B  (X   NNr�B  G?�      X   NNPr�B  G?�      uX   POSr�B  j�  �r�B  h h(h
c__builtin__
__main__
hNN}r�B  Ntr�B  Rr�B  �r�B  Rr�B  (X   VBZr�B  G?ٙ�����X   JJr�B  G?�333333uX   TOr�B  j)  �r�B  h h(h
c__builtin__
__main__
hNN}r�B  Ntr�B  Rr�B  �r�B  Rr�B  (X   VBr�B  G?��m��m�X   DTr�B  G?�I$�I$�X   WPr�B  G?�I$�I$�uX   PRPr�B  j�  �r�B  h h(h
c__builtin__
__main__
hNN}r�B  Ntr�B  Rr�B  �r�B  Rr�B  (X   JJr�B  G?ڪ�����X   NNr�B  G?�      X   INr�B  G?ʪ�����NG?�UUUUUUX   PRPr�B  G?�UUUUUUX   DTr�B  G?�UUUUUUuj�1  j�(  �r�B  h h(h
c__builtin__
__main__
hNN}r�B  Ntr�B  Rr�B  �r�B  Rr�B  (h�G?�I$�I$�X   INr�B  G?��m��m�X   DTr�B  G?�I$�I$�X   NNr�B  G?�m��m��uX   VBPr�B  j�  �r�B  h h(h
c__builtin__
__main__
hNN}r�B  Ntr�B  Rr�B  �r�B  Rr�B  (h�G?ٙ�����X   INr�B  G?ə�����X   NNPr�B  G?ə�����X   VBDr�B  G?ə�����uhMj�)  �r�B  h h(h
c__builtin__
__main__
hNN}r�B  Ntr�B  Rr�B  �r�B  Rr�B  (X   WPr�B  G?�wwwwwwX   WDTr�B  G?�UUUUUUX   CCr�B  G?�X   TOr�B  G?�X   NNr�B  G?�X   PRPr�B  G?�X   INr�B  G?�X   DTr�B  G?�uj�)  j�B  �r�B  h h(h
c__builtin__
__main__
hNN}r�B  Ntr�B  Rr�B  �r�B  Rr�B  (X   JJr�B  G?Ɩ�����X   VBPr�B  G?�X   VBZr�B  G?֖�����X   NNr�B  G?�X   VBDr�B  G?�X   MDr�B  G?�uh�j4  �r�B  h h(h
c__builtin__
__main__
hNN}r�B  Ntr�B  Rr�B  �r�B  Rr�B  (hMG?�E�t]FX   NNPr�B  G?�E�t]FX   JJr�B  G?�E�t]FX   WDTr�B  G?�t]E�tuj4  hM�r�B  h h(h
c__builtin__
__main__
hNN}r�B  Ntr�B  Rr�B  �r�B  Rr�B  (X   TOr C  G?�UUUUUUX   RBrC  G?�UUUUUUX   VBGrC  G?�UUUUUUuX   POSrC  j\  �rC  h h(h
c__builtin__
__main__
hNN}rC  NtrC  RrC  �rC  Rr	C  (X   MDr
C  G?�UUUUUUX   VBPrC  G?�UUUUUUuj)  j4  �rC  h h(h
c__builtin__
__main__
hNN}rC  NtrC  RrC  �rC  RrC  (X   NNrC  G?�      X   CDrC  G?�      X   NNSrC  G?�      h�G?�      uX   RBrC  j�*  �rC  h h(h
c__builtin__
__main__
hNN}rC  NtrC  RrC  �rC  RrC  (X   JJrC  G?�      X   INrC  G?�      X   VBNrC  G?�      uX   VBGrC  jH
  �r C  h h(h
c__builtin__
__main__
hNN}r!C  Ntr"C  Rr#C  �r$C  Rr%C  (X   NNSr&C  G?��!B�X   WPr'C  G?��!B�X   INr(C  G?��!B�X   WDTr)C  G?��!B�X   DTr*C  G?��1�c�X   JJr+C  G?��1�c�X   VBGr,C  G?��1�c�X   NNPr-C  G?��!B�X   PRPr.C  G?��!B�X   RBr/C  G?��!B�X   VBNr0C  G?��1�c�uX   RBSr1C  j^  �r2C  h h(h
c__builtin__
__main__
hNN}r3C  Ntr4C  Rr5C  �r6C  Rr7C  (X   DTr8C  G?���|X   NNr9C  G?�d�6M�eX   VBGr:C  G?�E�t]FX   PRP$r;C  G?�E�t]FX   JJr<C  G?�E�t]FX   VBNr=C  G?���|X   NNSr>C  G?�E�t]FX   WPr?C  G?���|X   CDr@C  G?���|h�G?���|uX   PRPrAC  jK$  �rBC  h h(h
c__builtin__
__main__
hNN}rCC  NtrDC  RrEC  �rFC  RrGC  (X   TOrHC  G?ٙ�����X   WRBrIC  G?�������X   INrJC  G?�333333X   JJrKC  G?�������h�G?�333333X   ''rLC  G?�������ujK$  jHC  �rMC  h h(h
c__builtin__
__main__
hNN}rNC  NtrOC  RrPC  �rQC  RrRC  (X   VBrSC  G?�|��|X   NNSrTC  G?���|X   DTrUC  G?�E�t]FX   TOrVC  G?���|X   JJSrWC  G?���|X   JJrXC  G?���|X   NNrYC  G?���|uX   JJRrZC  hM�r[C  h h(h
c__builtin__
__main__
hNN}r\C  Ntr]C  Rr^C  �r_C  Rr`C  (X   INraC  G?�333333X   NNPrbC  G?�333333X   JJRrcC  G?�333333X   DTrdC  G?�������X   oovreC  G?�������X   WPrfC  G?�333333X   VBNrgC  G?�������X   NNSrhC  G?�������uX   ''riC  j6  �rjC  h h(h
c__builtin__
__main__
hNN}rkC  NtrlC  RrmC  �rnC  RroC  (X   VBGrpC  G?�333333X   DTrqC  G?ٙ�����uX   NNPrrC  j�	  �rsC  h h(h
c__builtin__
__main__
hNN}rtC  NtruC  RrvC  �rwC  RrxC  (X   INryC  G?�!d,��X   NNrzC  G?��zoM�X   CCr{C  G?�B�Y!dX   JJr|C  G?��B�YX   TOr}C  G?�B�Y!dh�G?�B�Y!duj�
  j�  �r~C  h h(h
c__builtin__
__main__
hNN}rC  Ntr�C  Rr�C  �r�C  Rr�C  (X   JJr�C  G?�      h�G?�      X   PRP$r�C  G?�      uX   TOr�C  jP!  �r�C  h h(h
c__builtin__
__main__
hNN}r�C  Ntr�C  Rr�C  �r�C  Rr�C  (X   NNSr�C  G?؝�؝��X   INr�C  G?݉؝�؞X   JJr�C  G?ñ;�;uX   VBNr�C  jT#  �r�C  h h(h
c__builtin__
__main__
hNN}r�C  Ntr�C  Rr�C  �r�C  Rr�C  (X   RBr�C  G?�I$�I$�X   JJr�C  G?�I$�I$�X   RBSr�C  G?�I$�I$�uX   MDr�C  j�  �r�C  h h(h
c__builtin__
__main__
hNN}r�C  Ntr�C  Rr�C  �r�C  Rr�C  (X   NNSr�C  G?ñ;�;X   TOr�C  G?ñ;�;X   VBGr�C  G?ñ;�;X   DTr�C  G?͉؝�؞X   PRP$r�C  G?ñ;�;X   NNPr�C  G?ñ;�;uX   INr�C  N�r�C  h h(h
c__builtin__
__main__
hNN}r�C  Ntr�C  Rr�C  �r�C  Rr�C  NG?�      sX   TOr�C  j  �r�C  h h(h
c__builtin__
__main__
hNN}r�C  Ntr�C  Rr�C  �r�C  Rr�C  (X   INr�C  G?��m��m�X   NNr�C  G?�m��m��X   NNPr�C  G?�I$�I$�X   JJr�C  G?�I$�I$�X   NNSr�C  G?�I$�I$�uX   oovr�C  N�r�C  h h(h
c__builtin__
__main__
hNN}r�C  Ntr�C  Rr�C  �r�C  Rr�C  NG?�      sX   MDr�C  j�  �r�C  h h(h
c__builtin__
__main__
hNN}r�C  Ntr�C  Rr�C  �r�C  Rr�C  (X   INr�C  G?�      X   NNSr�C  G?�      uX   ''r�C  hM�r�C  h h(h
c__builtin__
__main__
hNN}r�C  Ntr�C  Rr�C  �r�C  Rr�C  (X   WRBr�C  G?�333333X   ``r�C  G?ə�����X   CCr�C  G?�333333X   WPr�C  G?�333333X   INr�C  G?�������X   NNPr�C  G?�������uX   VBZr�C  j�  �r�C  h h(h
c__builtin__
__main__
hNN}r�C  Ntr�C  Rr�C  �r�C  Rr�C  (X   VBNr�C  G?�����/hX   ''r�C  G?�q�q�h�G?�����/hX   NNSr�C  G?�����/hX   JJr�C  G?�����/hX   NNPr�C  G?�����/hX   VBr�C  G?�q�q�uj�
  j�C  �r�C  h h(h
c__builtin__
__main__
hNN}r�C  Ntr�C  Rr�C  �r�C  Rr�C  (X   NNr�C  G?�E�t]FX   VBNr�C  G?�E�t]FX   VBDr�C  G?�E�t]FX   VBZr�C  G?�E�t]FuX   WRBr�C  j�  �r�C  h h(h
c__builtin__
__main__
hNN}r�C  Ntr�C  Rr�C  �r�C  Rr�C  (X   VBPr�C  G?�I$�I$�X   VBDr�C  G?�m��m��X   JJr�C  G?�I$�I$�uh�j6  �r�C  h h(h
c__builtin__
__main__
hNN}r�C  Ntr�C  Rr�C  �r�C  Rr�C  X   VBDr�C  G?�      sX   WPr�C  j�#  �r D  h h(h
c__builtin__
__main__
hNN}rD  NtrD  RrD  �rD  RrD  (X   VBZrD  G?�I$�I$�X   MDrD  G?�I$�I$�X   VBDrD  G?�m��m��uX   WDTr	D  jk*  �r
D  h h(h
c__builtin__
__main__
hNN}rD  NtrD  RrD  �rD  RrD  (X   VBPrD  G?�m��m��X   VBDrD  G?�I$�I$�X   MDrD  G?�I$�I$�uX   WRBrD  j�  �rD  h h(h
c__builtin__
__main__
hNN}rD  NtrD  RrD  �rD  RrD  (X   NNSrD  G?�UUUUUUX   CCrD  G?�UUUUUUX   VBZrD  G?�UUUUUUuX   JJRrD  j 0  �rD  h h(h
c__builtin__
__main__
hNN}rD  Ntr D  Rr!D  �r"D  Rr#D  (h�G?�333333X   NNSr$D  G?ə�����X   INr%D  G?ə�����uX   RPr&D  j�,  �r'D  h h(h
c__builtin__
__main__
hNN}r(D  Ntr)D  Rr*D  �r+D  Rr,D  (X   VBZr-D  G?�E�t]FX   INr.D  G?�E�t]h�G?�E�t]FX   DTr/D  G?�E�t]FuX   ''r0D  j�  �r1D  h h(h
c__builtin__
__main__
hNN}r2D  Ntr3D  Rr4D  �r5D  Rr6D  (X   VBDr7D  G?�      h�G?�      X   DTr8D  G?�      uX   oovr9D  j0  �r:D  h h(h
c__builtin__
__main__
hNN}r;D  Ntr<D  Rr=D  �r>D  Rr?D  (X   oovr@D  G?�X   VBPrAD  G?�X   MDrBD  G?ə�����X   INrCD  G?�X   RBrDD  G?�uj�9  j�=  �rED  h h(h
c__builtin__
__main__
hNN}rFD  NtrGD  RrHD  �rID  RrJD  (X   VBDrKD  G?�      X   VBPrLD  G?�      uX   DTrMD  j�  �rND  h h(h
c__builtin__
__main__
hNN}rOD  NtrPD  RrQD  �rRD  RrSD  (X   NNPrTD  G?ñ;�;X   VBrUD  G?�'bv'bvX   JJrVD  G?ñ;�;uX   VBGrWD  j�'  �rXD  h h(h
c__builtin__
__main__
hNN}rYD  NtrZD  Rr[D  �r\D  Rr]D  (X   WRBr^D  G?�E�t]FX   TOr_D  G?�E�t]FX   INr`D  G?�t]E�th�G?�E�t]FX   NNraD  G?�E�t]FuX   ''rbD  j�  �rcD  h h(h
c__builtin__
__main__
hNN}rdD  NtreD  RrfD  �rgD  RrhD  (X   NNriD  G?�333333X   VBZrjD  G?ٙ�����uji)  j�:  �rkD  h h(h
c__builtin__
__main__
hNN}rlD  NtrmD  RrnD  �roD  RrpD  (X   oovrqD  G?�333333X   CCrrD  G?ٙ�����uj�:  jqD  �rsD  h h(h
c__builtin__
__main__
hNN}rtD  NtruD  RrvD  �rwD  RrxD  (X   CCryD  G?�UUUUUUX   VBGrzD  G?�q�q�X   VBNr{D  G?�q�q�X   DTr|D  G?�q�q�uj  j�9  �r}D  h h(h
c__builtin__
__main__
hNN}r~D  NtrD  Rr�D  �r�D  Rr�D  (X   INr�D  G?�I$�I$�X   DTr�D  G?�m��m��X   RBr�D  G?�I$�I$�uX   VBGr�D  j�	  �r�D  h h(h
c__builtin__
__main__
hNN}r�D  Ntr�D  Rr�D  �r�D  Rr�D  (X   TOr�D  G?�      X   INr�D  G?�      uX   WRBr�D  hM�r�D  h h(h
c__builtin__
__main__
hNN}r�D  Ntr�D  Rr�D  �r�D  Rr�D  (X   INr�D  G?�      X   JJr�D  G?�UUUUUUX   CCr�D  G?�UUUUUUX   RBr�D  G?�UUUUUUuX   VBPr�D  N�r�D  h h(h
c__builtin__
__main__
hNN}r�D  Ntr�D  Rr�D  �r�D  Rr�D  NG?�      sX   WRBr�D  j�  �r�D  h h(h
c__builtin__
__main__
hNN}r�D  Ntr�D  Rr�D  �r�D  Rr�D  (X   NNPr�D  G?�      X   NNr�D  G?�      uNh5�r�D  h h(h
c__builtin__
__main__
hNN}r�D  Ntr�D  Rr�D  �r�D  Rr�D  (X   NNSr�D  G?�E�t]FX   PRPr�D  G?�E�t]FX   WPr�D  G?�E�t]FX   PRP$r�D  G?�E�t]FX   oovr�D  G?�t]E�tujFA  j20  �r�D  h h(h
c__builtin__
__main__
hNN}r�D  Ntr�D  Rr�D  �r�D  Rr�D  (X   VBr�D  G?�q�q�X   WDTr�D  G?�q�q�X   DTr�D  G?�UUUUUUuX   MDr�D  j
"  �r�D  h h(h
c__builtin__
__main__
hNN}r�D  Ntr�D  Rr�D  �r�D  Rr�D  (X   NNr�D  G?��q�rX   VBGr�D  G?�q�q�X   JJr�D  G?�q�q�uh�j7  �r�D  h h(h
c__builtin__
__main__
hNN}r�D  Ntr�D  Rr�D  �r�D  Rr�D  (X   VBZr�D  G?�UUUUUUX   JJr�D  G?�UUUUUUX   VBPr�D  G?�UUUUUUuX   MDr�D  j�  �r�D  h h(h
c__builtin__
__main__
hNN}r�D  Ntr�D  Rr�D  �r�D  Rr�D  (X   NNSr�D  G?�333333X   INr�D  G?ٙ�����uX   TOr�D  j�  �r�D  h h(h
c__builtin__
__main__
hNN}r�D  Ntr�D  Rr�D  �r�D  Rr�D  (X   JJr�D  G?��m��m�X   RBr�D  G?�I$�I$�uX   NNr�D  j(  �r�D  h h(h
c__builtin__
__main__
hNN}r�D  Ntr�D  Rr�D  �r�D  Rr�D  (X   NNSr�D  G?Ǵ%�	{BX   VBPr�D  G?�����/hX   NNr�D  G?Ǵ%�	{BX   RBr�D  G?�����/hX   TOr�D  G?�q�q�X   INr�D  G?�q�q�X   VBNr�D  G?�����/hX   JJr�D  G?�����/hujz  j6/  �r�D  h h(h
c__builtin__
__main__
hNN}r�D  Ntr�D  Rr�D  �r�D  Rr�D  (X   NNPr�D  G?�E�t]FX   NNr�D  G?�E�t]FX   NNSr�D  G?�E�t]FX   JJr�D  G?�t]E�tuX   PRPr�D  j�  �r�D  h h(h
c__builtin__
__main__
hNN}r�D  Ntr�D  Rr E  �rE  RrE  (X   NNrE  G?�      X   JJrE  G?�      uX   JJRrE  jIC  �rE  h h(h
c__builtin__
__main__
hNN}rE  NtrE  Rr	E  �r
E  RrE  X   PRPrE  G?�      sX   JJRrE  j0  �rE  h h(h
c__builtin__
__main__
hNN}rE  NtrE  RrE  �rE  RrE  (X   NNrE  G?͉؝�؞X   NNSrE  G?݉؝�؞X   DTrE  G?ӱ;�;uX   oovrE  j�>  �rE  h h(h
c__builtin__
__main__
hNN}rE  NtrE  RrE  �rE  RrE  (X   NNrE  G?�I$�I$�X   JJrE  G?�I$�I$�X   PRPr E  G?�m��m��uX   RBr!E  jt#  �r"E  h h(h
c__builtin__
__main__
hNN}r#E  Ntr$E  Rr%E  �r&E  Rr'E  (X   JJr(E  G?�      X   RBr)E  G?�      X   DTr*E  G?�      h�G?�      X   NNPr+E  G?�      X   INr,E  G?�      uX   JJSr-E  jT  �r.E  h h(h
c__builtin__
__main__
hNN}r/E  Ntr0E  Rr1E  �r2E  Rr3E  (X   NNr4E  G?͉؝�؞X   CDr5E  G?ñ;�;X   WPr6E  G?ñ;�;X   VBPr7E  G?݉؝�؞uj$
  j�/  �r8E  h h(h
c__builtin__
__main__
hNN}r9E  Ntr:E  Rr;E  �r<E  Rr=E  (X   RBr>E  G?�X   DTr?E  G?�X   NNr@E  G?�h�G?�hMG?�X   NNSrAE  G?�X   CDrBE  G?ə�����uX   WPrCE  jz  �rDE  h h(h
c__builtin__
__main__
hNN}rEE  NtrFE  RrGE  �rHE  RrIE  (X   WPrJE  G?�UUUUUUX   WRBrKE  G?�UUUUUUX   RBrLE  G?�UUUUUUuX   WDTrME  jR*  �rNE  h h(h
c__builtin__
__main__
hNN}rOE  NtrPE  RrQE  �rRE  RrSE  X   NNrTE  G?�      sX   MDrUE  jU  �rVE  h h(h
c__builtin__
__main__
hNN}rWE  NtrXE  RrYE  �rZE  Rr[E  (X   VBr\E  G?�      X   DTr]E  G?�      uX   VBNr^E  j@  �r_E  h h(h
c__builtin__
__main__
hNN}r`E  NtraE  RrbE  �rcE  RrdE  X   VBreE  G?�      sX   ``rfE  j  �rgE  h h(h
c__builtin__
__main__
hNN}rhE  NtriE  RrjE  �rkE  RrlE  (X   PRPrmE  G?�I$�I$�X   ''rnE  G?�I$�I$�X   ``roE  G?�m��m��uh�j�  �rpE  h h(h
c__builtin__
__main__
hNN}rqE  NtrrE  RrsE  �rtE  RruE  (h�G?�m��m��X   CCrvE  G?�I$�I$�NG?�I$�I$�uX   WDTrwE  j9  �rxE  h h(h
c__builtin__
__main__
hNN}ryE  NtrzE  Rr{E  �r|E  Rr}E  (X   JJr~E  G?�      h�G?�      uX   TOrE  j  �r�E  h h(h
c__builtin__
__main__
hNN}r�E  Ntr�E  Rr�E  �r�E  Rr�E  (X   NNr�E  G?�B�Y!dX   NNSr�E  G?�B�Y!dX   CCr�E  G?�B�Y!dX   VBGr�E  G?�B�Y!dX   VBr�E  G?��B�YX   JJr�E  G?�B�Y!dX   ``r�E  G?�B�Y!duX   WPr�E  j  �r�E  h h(h
c__builtin__
__main__
hNN}r�E  Ntr�E  Rr�E  �r�E  Rr�E  (X   INr�E  G?�      X   JJr�E  G?�      X   NNPr�E  G?�      X   PRP$r�E  G?�      X   TOr�E  G?�      uj5  jQ  �r�E  h h(h
c__builtin__
__main__
hNN}r�E  Ntr�E  Rr�E  �r�E  Rr�E  (X   VBr�E  G?�      X   NNPr�E  G?�      X   DTr�E  G?�      uX   POSr�E  j`  �r�E  h h(h
c__builtin__
__main__
hNN}r�E  Ntr�E  Rr�E  �r�E  Rr�E  X   NNSr�E  G?�      sj 1  hM�r�E  h h(h
c__builtin__
__main__
hNN}r�E  Ntr�E  Rr�E  �r�E  Rr�E  (X   CCr�E  G?ə�����X   DTr�E  G?ə�����X   WPr�E  G?ə�����X   WDTr�E  G?�X   VBGr�E  G?�X   WRBr�E  G?�uX   VBPr�E  j�7  �r�E  h h(h
c__builtin__
__main__
hNN}r�E  Ntr�E  Rr�E  �r�E  Rr�E  (X   VBNr�E  G?�X   NNr�E  G?�X   NNSr�E  G?�X   JJr�E  G?ə�����X   VBDr�E  G?�X   NNPr�E  G?�uX   JJRr�E  j+7  �r�E  h h(h
c__builtin__
__main__
hNN}r�E  Ntr�E  Rr�E  �r�E  Rr�E  (X   NNr�E  G?�m��m��X   VBNr�E  G?�I$�I$�X   CDr�E  G?�I$�I$�uX   MDr�E  j"  �r�E  h h(h
c__builtin__
__main__
hNN}r�E  Ntr�E  Rr�E  �r�E  Rr�E  X   JJr�E  G?�      sX   VBr�E  j7  �r�E  h h(h
c__builtin__
__main__
hNN}r�E  Ntr�E  Rr�E  �r�E  Rr�E  (X   JJr�E  G?�X   RBr�E  G?Ɩ�����X   NNSr�E  G?�h�G?�X   NNr�E  G?�X   INr�E  G?�ujC  j�)  �r�E  h h(h
c__builtin__
__main__
hNN}r�E  Ntr�E  Rr�E  �r�E  Rr�E  (X   VBDr�E  G?ڪ�����X   VBZr�E  G?�UUUUUUX   MDr�E  G?�UUUUUUX   VBPr�E  G?�      uj�  jYB  �r�E  h h(h
c__builtin__
__main__
hNN}r�E  Ntr�E  Rr�E  �r�E  Rr�E  X   VBZr�E  G?�      sX   POSr�E  ja  �r�E  h h(h
c__builtin__
__main__
hNN}r�E  Ntr�E  Rr�E  �r�E  Rr�E  (h�G?�      X   NNr�E  G?�      X   RPr�E  G?�      X   INr�E  G?�      X   NNPr�E  G?�      X   DTr�E  G?�      ujQ  hM�r�E  h h(h
c__builtin__
__main__
hNN}r�E  Ntr F  RrF  �rF  RrF  (X   WPrF  G?�q�q�X   WRBrF  G?�q�q�X   CCrF  G?�q�q�X   oovrF  G?�q�q�X   VBDrF  G?�q�q�X   NNr	F  G?�q�q�X   DTr
F  G?�q�q�X   ``rF  G?�q�q�uX   PRPrF  j�0  �rF  h h(h
c__builtin__
__main__
hNN}rF  NtrF  RrF  �rF  RrF  (h�G?�      X   NNrF  G?�      X   NNSrF  G?�      X   INrF  G?�      X   VBZrF  G?�      X   PRPrF  G?�      uj�.  j�-  �rF  h h(h
c__builtin__
__main__
hNN}rF  NtrF  RrF  �rF  RrF  (X   NNPrF  G?�q�q�X   NNrF  G?�UUUUUUX   NNSr F  G?�q�q�h�G?�q�q�uX   JJRr!F  jb  �r"F  h h(h
c__builtin__
__main__
hNN}r#F  Ntr$F  Rr%F  �r&F  Rr'F  (X   NNSr(F  G?�E�t]h�G?�E�t]FX   INr)F  G?�      X   JJr*F  G?�E�t]FX   VBNr+F  G?�E�t]FuX   oovr,F  jIA  �r-F  h h(h
c__builtin__
__main__
hNN}r.F  Ntr/F  Rr0F  �r1F  Rr2F  (X   NNr3F  G?�      NG?�      h�G?�      X   VBNr4F  G?�      uX   RBSr5F  j�8  �r6F  h h(h
c__builtin__
__main__
hNN}r7F  Ntr8F  Rr9F  �r:F  Rr;F  X   NNr<F  G?�      sX   VBGr=F  N�r>F  h h(h
c__builtin__
__main__
hNN}r?F  Ntr@F  RrAF  �rBF  RrCF  NG?�      sX   WDTrDF  j:  �rEF  h h(h
c__builtin__
__main__
hNN}rFF  NtrGF  RrHF  �rIF  RrJF  (X   INrKF  G?�      X   VBDrLF  G?�      uX   JJrMF  N�rNF  h h(h
c__builtin__
__main__
hNN}rOF  NtrPF  RrQF  �rRF  RrSF  NG?�      sX   POSrTF  jb  �rUF  h h(h
c__builtin__
__main__
hNN}rVF  NtrWF  RrXF  �rYF  RrZF  (X   RBr[F  G?ٙ�����X   VBr\F  G?�333333uX   INr]F  j�  �r^F  h h(h
c__builtin__
__main__
hNN}r_F  Ntr`F  RraF  �rbF  RrcF  X   NNrdF  G?�      sX   PRP$reF  j�  �rfF  h h(h
c__builtin__
__main__
hNN}rgF  NtrhF  RriF  �rjF  RrkF  (X   DTrlF  G?�      hMG?�      uX   NNSrmF  j�  �rnF  h h(h
c__builtin__
__main__
hNN}roF  NtrpF  RrqF  �rrF  RrsF  (X   VBPrtF  G?�UUUUUUX   INruF  G?�UUUUUUX   CCrvF  G?�UUUUUUuj�  j30  �rwF  h h(h
c__builtin__
__main__
hNN}rxF  NtryF  RrzF  �r{F  Rr|F  (X   NNSr}F  G?�B�Y!dX   NNPr~F  G?вB�YX   RPrF  G?�B�Y!dX   INr�F  G?��B�Yh�G?�B�Y!dX   NNr�F  G?�B�Y!dX   TOr�F  G?�B�Y!dX   DTr�F  G?�B�Y!duh�j�  �r�F  h h(h
c__builtin__
__main__
hNN}r�F  Ntr�F  Rr�F  �r�F  Rr�F  X   PRPr�F  G?�      sX   WDTr�F  j�  �r�F  h h(h
c__builtin__
__main__
hNN}r�F  Ntr�F  Rr�F  �r�F  Rr�F  X   VBDr�F  G?�      sX   RBr�F  jq  �r�F  h h(h
c__builtin__
__main__
hNN}r�F  Ntr�F  Rr�F  �r�F  Rr�F  (X   VBPr�F  G?��m��m�X   VBDr�F  G?�I$�I$�uji:  j�1  �r�F  h h(h
c__builtin__
__main__
hNN}r�F  Ntr�F  Rr�F  �r�F  Rr�F  X   NNr�F  G?�      sNh6�r�F  h h(h
c__builtin__
__main__
hNN}r�F  Ntr�F  Rr�F  �r�F  Rr�F  X   INr�F  G?�      sX   MDr�F  j�  �r�F  h h(h
c__builtin__
__main__
hNN}r�F  Ntr�F  Rr�F  �r�F  Rr�F  X   WPr�F  G?�      sX   VBr�F  j.  �r�F  h h(h
c__builtin__
__main__
hNN}r�F  Ntr�F  Rr�F  �r�F  Rr�F  (X   TOr�F  G?Ɩ�����X   INr�F  G?�X   VBr�F  G?�h�G?�X   RBr�F  G?�X   CDr�F  G?�uX   RPr�F  j�$  �r�F  h h(h
c__builtin__
__main__
hNN}r�F  Ntr�F  Rr�F  �r�F  Rr�F  (X   INr�F  G?�      X   NNr�F  G?�      X   NNSr�F  G?�      uX   RBSr�F  j�8  �r�F  h h(h
c__builtin__
__main__
hNN}r�F  Ntr�F  Rr�F  �r�F  Rr�F  (X   VBNr�F  G?�UUUUUUX   INr�F  G?�UUUUUUh�G?�UUUUUUuX   JJRr�F  j0  �r�F  h h(h
c__builtin__
__main__
hNN}r�F  Ntr�F  Rr�F  �r�F  Rr�F  X   INr�F  G?�      sX   JJRr�F  jn?  �r�F  h h(h
c__builtin__
__main__
hNN}r�F  Ntr�F  Rr�F  �r�F  Rr�F  X   RBr�F  G?�      sX   MDr�F  j"  �r�F  h h(h
c__builtin__
__main__
hNN}r�F  Ntr�F  Rr�F  �r�F  Rr�F  X   VBr�F  G?�      sX   POSr�F  j  �r�F  h h(h
c__builtin__
__main__
hNN}r�F  Ntr�F  Rr�F  �r�F  Rr�F  X   DTr�F  G?�      shMj�9  �r�F  h h(h
c__builtin__
__main__
hNN}r�F  Ntr�F  Rr�F  �r�F  Rr�F  X   JJr�F  G?�      sj�@  N�r�F  h h(h
c__builtin__
__main__
hNN}r�F  Ntr�F  Rr�F  �r�F  Rr�F  NG?�      sj�?  N�r�F  h h(h
c__builtin__
__main__
hNN}r�F  Ntr G  RrG  �rG  RrG  NG?�      sX   VBDrG  N�rG  h h(h
c__builtin__
__main__
hNN}rG  NtrG  RrG  �r	G  Rr
G  NG?�      sX   WPrG  N�rG  h h(h
c__builtin__
__main__
hNN}rG  NtrG  RrG  �rG  RrG  NG?�      sX   VBZrG  N�rG  h h(h
c__builtin__
__main__
hNN}rG  NtrG  RrG  �rG  RrG  NG?�      sX   WRBrG  N�rG  h h(h
c__builtin__
__main__
hNN}rG  NtrG  RrG  �rG  RrG  NG?�      sX   CCr G  N�r!G  h h(h
c__builtin__
__main__
hNN}r"G  Ntr#G  Rr$G  �r%G  Rr&G  NG?�      sX   ''r'G  j�B  �r(G  h h(h
c__builtin__
__main__
hNN}r)G  Ntr*G  Rr+G  �r,G  Rr-G  X   MDr.G  G?�      sX   NNPSr/G  j3  �r0G  h h(h
c__builtin__
__main__
hNN}r1G  Ntr2G  Rr3G  �r4G  Rr5G  (X   NNr6G  G?؝�؝��X   JJr7G  G?ñ;�;X   VBNr8G  G?ñ;�;h�G?ӱ;�;uj�<  jnE  �r9G  h h(h
c__builtin__
__main__
hNN}r:G  Ntr;G  Rr<G  �r=G  Rr>G  X   VBr?G  G?�      sj�  jL<  �r@G  h h(h
c__builtin__
__main__
hNN}rAG  NtrBG  RrCG  �rDG  RrEG  (h�G?�UUUUUUX   NNrFG  G?�UUUUUUuX   RBSrGG  j�C  �rHG  h h(h
c__builtin__
__main__
hNN}rIG  NtrJG  RrKG  �rLG  RrMG  X   JJrNG  G?�      sX   TOrOG  hM�rPG  h h(h
c__builtin__
__main__
hNN}rQG  NtrRG  RrSG  �rTG  RrUG  (X   VBGrVG  G?�q�q�X   RBrWG  G?�q�q�X   INrXG  G?�UUUUUUX   TOrYG  G?�q�q�uX   DTrZG  j�  �r[G  h h(h
c__builtin__
__main__
hNN}r\G  Ntr]G  Rr^G  �r_G  Rr`G  (X   JJraG  G?�m��m��X   DTrbG  G?�I$�I$�X   VBZrcG  G?�I$�I$�uX   NNPSrdG  j3  �reG  h h(h
c__builtin__
__main__
hNN}rfG  NtrgG  RrhG  �riG  RrjG  (h�G?�UUUUUUX   PRPrkG  G?�UUUUUUX   DTrlG  G?�UUUUUUuX   CCrmG  h��rnG  h h(h
c__builtin__
__main__
hNN}roG  NtrpG  RrqG  �rrG  RrsG  NG?�      sh�j�  �rtG  h h(h
c__builtin__
__main__
hNN}ruG  NtrvG  RrwG  �rxG  RryG  (X   NNPrzG  G?�      X   NNr{G  G?�      X   JJr|G  G?�      uX   INr}G  j\  �r~G  h h(h
c__builtin__
__main__
hNN}rG  Ntr�G  Rr�G  �r�G  Rr�G  X   DTr�G  G?�      shMhM�r�G  h h(h
c__builtin__
__main__
hNN}r�G  Ntr�G  Rr�G  �r�G  Rr�G  (X   WRBr�G  G?�      X   NNr�G  G?�      uX   ''r�G  j=  �r�G  h h(h
c__builtin__
__main__
hNN}r�G  Ntr�G  Rr�G  �r�G  Rr�G  X   RBr�G  G?�      sh�j;  �r�G  h h(h
c__builtin__
__main__
hNN}r�G  Ntr�G  Rr�G  �r�G  Rr�G  X   NNPr�G  G?�      sj>  jjD  �r�G  h h(h
c__builtin__
__main__
hNN}r�G  Ntr�G  Rr�G  �r�G  Rr�G  (X   INr�G  G?�������X   RPr�G  G?�������X   JJr�G  G?�������X   VBr�G  G?�������X   DTr�G  G?ə�����X   PRP$r�G  G?�������X   ``r�G  G?�������X   VBNr�G  G?�������X   NNSr�G  G?�������uX   TOr�G  N�r�G  h h(h
c__builtin__
__main__
hNN}r�G  Ntr�G  Rr�G  �r�G  Rr�G  NG?�      sX   POSr�G  N�r�G  h h(h
c__builtin__
__main__
hNN}r�G  Ntr�G  Rr�G  �r�G  Rr�G  NG?�      sX   RBSr�G  N�r�G  h h(h
c__builtin__
__main__
hNN}r�G  Ntr�G  Rr�G  �r�G  Rr�G  NG?�      sX   PRPr�G  N�r�G  h h(h
c__builtin__
__main__
hNN}r�G  Ntr�G  Rr�G  �r�G  Rr�G  NG?�      sX   CCr�G  j�  �r�G  h h(h
c__builtin__
__main__
hNN}r�G  Ntr�G  Rr�G  �r�G  Rr�G  (X   NNr�G  G?�      X   DTr�G  G?�      X   NNSr�G  G?�      X   JJr�G  G?�      X   PRP$r�G  G?�      X   oovr�G  G?�      X   VBr�G  G?�      uX   RBr�G  jE(  �r�G  h h(h
c__builtin__
__main__
hNN}r�G  Ntr�G  Rr�G  �r�G  Rr�G  (X   JJr�G  G?�UUUUUUX   NNr�G  G?�q�q�X   NNSr�G  G?�q�q�uX   JJSr�G  j�  �r�G  h h(h
c__builtin__
__main__
hNN}r�G  Ntr�G  Rr�G  �r�G  Rr�G  (X   VBPr�G  G?�      X   INr�G  G?�      uh�hM�r�G  h h(h
c__builtin__
__main__
hNN}r�G  Ntr�G  Rr�G  �r�G  Rr�G  (X   NNPr�G  G?�      h�G?�      uX   PRP$r�G  hM�r�G  h h(h
c__builtin__
__main__
hNN}r�G  Ntr�G  Rr�G  �r�G  Rr�G  X   WPr�G  G?�      sX   POSr�G  jc  �r�G  h h(h
c__builtin__
__main__
hNN}r�G  Ntr�G  Rr�G  �r�G  Rr�G  (X   NNr�G  G?�UUUUUUX   MDr�G  G?�UUUUUUX   VBDr H  G?�UUUUUUuX   RPrH  N�rH  h h(h
c__builtin__
__main__
hNN}rH  NtrH  RrH  �rH  RrH  NG?�      sh�j<  �rH  h h(h
c__builtin__
__main__
hNN}r	H  Ntr
H  RrH  �rH  RrH  X   VBGrH  G?�      sX   oovrH  j�  �rH  h h(h
c__builtin__
__main__
hNN}rH  NtrH  RrH  �rH  RrH  X   INrH  G?�      sX   PRP$rH  j�  �rH  h h(h
c__builtin__
__main__
hNN}rH  NtrH  RrH  �rH  RrH  (X   JJrH  G?�333333X   NNrH  G?ٙ�����ujE  j.  �r H  h h(h
c__builtin__
__main__
hNN}r!H  Ntr"H  Rr#H  �r$H  Rr%H  X   RBr&H  G?�      sX   ``r'H  j�  �r(H  h h(h
c__builtin__
__main__
hNN}r)H  Ntr*H  Rr+H  �r,H  Rr-H  (X   PRPr.H  G?�I$�I$�X   VBZr/H  G?�I$�I$�X   VBr0H  G?�I$�I$�X   VBDr1H  G?�I$�I$�X   DTr2H  G?�I$�I$�X   NNSr3H  G?�I$�I$�uX   JJRr4H  jLC  �r5H  h h(h
c__builtin__
__main__
hNN}r6H  Ntr7H  Rr8H  �r9H  Rr:H  (X   VBr;H  G?�      X   NNr<H  G?�      uX   RBSr=H  j)9  �r>H  h h(h
c__builtin__
__main__
hNN}r?H  Ntr@H  RrAH  �rBH  RrCH  X   NNrDH  G?�      su(X   VBNrEH  j�  �rFH  h h(h
c__builtin__
__main__
hNN}rGH  NtrHH  RrIH  �rJH  RrKH  (X   WDTrLH  G?�UUUUUUh�G?�UUUUUUX   VBNrMH  G?�UUUUUUuX   WRBrNH  j�  �rOH  h h(h
c__builtin__
__main__
hNN}rPH  NtrQH  RrRH  �rSH  RrTH  (X   INrUH  G?�      X   NNSrVH  G?�      uj�  N�rWH  h h(h
c__builtin__
__main__
hNN}rXH  NtrYH  RrZH  �r[H  Rr\H  NG?�      sX   RPr]H  j%  �r^H  h h(h
c__builtin__
__main__
hNN}r_H  Ntr`H  RraH  �rbH  RrcH  (X   INrdH  G?�      X   NNPreH  G?�      X   TOrfH  G?�      h�G?�      uX   RBSrgH  j_  �rhH  h h(h
c__builtin__
__main__
hNN}riH  NtrjH  RrkH  �rlH  RrmH  h�G?�      sX   CCrnH  j�  �roH  h h(h
c__builtin__
__main__
hNN}rpH  NtrqH  RrrH  �rsH  RrtH  (X   ''ruH  G?�      X   NNPrvH  G?�      uX   RPrwH  je;  �rxH  h h(h
c__builtin__
__main__
hNN}ryH  NtrzH  Rr{H  �r|H  Rr}H  h�G?�      sX   MDr~H  jN@  �rH  h h(h
c__builtin__
__main__
hNN}r�H  Ntr�H  Rr�H  �r�H  Rr�H  (X   DTr�H  G?�      X   VBr�H  G?�      uX   PRPr�H  jd   �r�H  h h(h
c__builtin__
__main__
hNN}r�H  Ntr�H  Rr�H  �r�H  Rr�H  X   JJr�H  G?�      sX   PRPr�H  j  �r�H  h h(h
c__builtin__
__main__
hNN}r�H  Ntr�H  Rr�H  �r�H  Rr�H  (X   JJr�H  G?�UUUUUUX   VBPr�H  G?�UUUUUUh�G?�UUUUUUuX   ``r�H  j�  �r�H  h h(h
c__builtin__
__main__
hNN}r�H  Ntr�H  Rr�H  �r�H  Rr�H  (X   VBPr�H  G?ٙ�����X   ''r�H  G?�333333uX   MDr�H  jF*  �r�H  h h(h
c__builtin__
__main__
hNN}r�H  Ntr�H  Rr�H  �r�H  Rr�H  h�G?�      sX   JJSr�H  j|%  �r�H  h h(h
c__builtin__
__main__
hNN}r�H  Ntr�H  Rr�H  �r�H  Rr�H  X   NNr�H  G?�      sX   VBZr�H  j�
  �r�H  h h(h
c__builtin__
__main__
hNN}r�H  Ntr�H  Rr�H  �r�H  Rr�H  (X   DTr�H  G?�      X   NNr�H  G?�      uX   RPr�H  j  �r�H  h h(h
c__builtin__
__main__
hNN}r�H  Ntr�H  Rr�H  �r�H  Rr�H  (X   VBZr�H  G?�      h�G?�      uX   CDr�H  jE  �r�H  h h(h
c__builtin__
__main__
hNN}r�H  Ntr�H  Rr�H  �r�H  Rr�H  X   CDr�H  G?�      sX   VBDr�H  j�  �r�H  h h(h
c__builtin__
__main__
hNN}r�H  Ntr�H  Rr�H  �r�H  Rr�H  (X   JJr�H  G?�UUUUUUX   ''r�H  G?ڪ�����X   NNPr�H  G?�      X   NNr�H  G?�UUUUUUujW  j2  �r�H  h h(h
c__builtin__
__main__
hNN}r�H  Ntr�H  Rr�H  �r�H  Rr�H  X   VBr�H  G?�      sX   ``r�H  j�  �r�H  h h(h
c__builtin__
__main__
hNN}r�H  Ntr�H  Rr�H  �r�H  Rr�H  (X   JJr�H  G?�      X   ''r�H  G?�      X   DTr�H  G?�      X   NNSr�H  G?�      X   VBNr�H  G?�      X   VBZr�H  G?�      X   VBr�H  G?�      uX   oovr�H  j#0  �r�H  h h(h
c__builtin__
__main__
hNN}r�H  Ntr�H  Rr�H  �r�H  Rr�H  X   NNr�H  G?�      sX   WDTr�H  j<  �r�H  h h(h
c__builtin__
__main__
hNN}r�H  Ntr�H  Rr�H  �r�H  Rr�H  h�G?�      sX   ''r�H  j�  �r�H  h h(h
c__builtin__
__main__
hNN}r�H  Ntr�H  Rr�H  �r�H  Rr�H  NG?�      sh�j�  �r�H  h h(h
c__builtin__
__main__
hNN}r I  NtrI  RrI  �rI  RrI  X   NNrI  G?�      sX   RPrI  j	4  �rI  h h(h
c__builtin__
__main__
hNN}rI  Ntr	I  Rr
I  �rI  RrI  X   NNPrI  G?�      shMh��rI  h h(h
c__builtin__
__main__
hNN}rI  NtrI  RrI  �rI  RrI  NG?�      sX   WRBrI  j�-  �rI  h h(h
c__builtin__
__main__
hNN}rI  NtrI  RrI  �rI  RrI  h�G?�      shMN�rI  h h(h
c__builtin__
__main__
hNN}rI  NtrI  RrI  �rI  Rr I  NG?�      sX   MDr!I  j�  �r"I  h h(h
c__builtin__
__main__
hNN}r#I  Ntr$I  Rr%I  �r&I  Rr'I  (X   JJr(I  G?�      X   NNSr)I  G?�      uX   DTr*I  N�r+I  h h(h
c__builtin__
__main__
hNN}r,I  Ntr-I  Rr.I  �r/I  Rr0I  NG?�      sX   POSr1I  jd  �r2I  h h(h
c__builtin__
__main__
hNN}r3I  Ntr4I  Rr5I  �r6I  Rr7I  X   NNr8I  G?�      sh�j?  �r9I  h h(h
c__builtin__
__main__
hNN}r:I  Ntr;I  Rr<I  �r=I  Rr>I  (X   MDr?I  G?ٙ�����X   VBZr@I  G?�333333uX   WPrAI  j  �rBI  h h(h
c__builtin__
__main__
hNN}rCI  NtrDI  RrEI  �rFI  RrGI  (X   VBDrHI  G?�      X   VBPrII  G?�      uX   WPrJI  j  �rKI  h h(h
c__builtin__
__main__
hNN}rLI  NtrMI  RrNI  �rOI  RrPI  X   JJrQI  G?�      sX   RBSrRI  j4  �rSI  h h(h
c__builtin__
__main__
hNN}rTI  NtrUI  RrVI  �rWI  RrXI  (X   DTrYI  G?ٙ�����X   INrZI  G?�333333uj�  j1  �r[I  h h(h
c__builtin__
__main__
hNN}r\I  Ntr]I  Rr^I  �r_I  Rr`I  (X   VBraI  G?�333333X   MDrbI  G?ٙ�����uX   JJSrcI  j�?  �rdI  h h(h
c__builtin__
__main__
hNN}reI  NtrfI  RrgI  �rhI  RriI  h�G?�      sX   WDTrjI  j�  �rkI  h h(h
c__builtin__
__main__
hNN}rlI  NtrmI  RrnI  �roI  RrpI  X   VBZrqI  G?�      sX   RBSrrI  jI:  �rsI  h h(h
c__builtin__
__main__
hNN}rtI  NtruI  RrvI  �rwI  RrxI  X   NNryI  G?�      sj2&  hM�rzI  h h(h
c__builtin__
__main__
hNN}r{I  Ntr|I  Rr}I  �r~I  RrI  X   WPr�I  G?�      sX   RPr�I  j4  �r�I  h h(h
c__builtin__
__main__
hNN}r�I  Ntr�I  Rr�I  �r�I  Rr�I  X   DTr�I  G?�      sj�  j�6  �r�I  h h(h
c__builtin__
__main__
hNN}r�I  Ntr�I  Rr�I  �r�I  Rr�I  (X   ``r�I  G?�I$�I$�X   PRPr�I  G?�I$�I$�X   DTr�I  G?�I$�I$�X   RBr�I  G?�I$�I$�X   VBDr�I  G?�I$�I$�X   WRBr�I  G?�I$�I$�uX   ``r�I  N�r�I  h h(h
c__builtin__
__main__
hNN}r�I  Ntr�I  Rr�I  �r�I  Rr�I  NG?�      sh�j�  �r�I  h h(h
c__builtin__
__main__
hNN}r�I  Ntr�I  Rr�I  �r�I  Rr�I  X   NNPr�I  G?�      sj�&  j`B  �r�I  h h(h
c__builtin__
__main__
hNN}r�I  Ntr�I  Rr�I  �r�I  Rr�I  (X   JJr�I  G?�333333X   NNr�I  G?ٙ�����uX   ``r�I  j  �r�I  h h(h
c__builtin__
__main__
hNN}r�I  Ntr�I  Rr�I  �r�I  Rr�I  (X   VBZr�I  G?�333333X   JJr�I  G?�333333X   NNr�I  G?ə�����X   VBDr�I  G?ə�����uX   JJRr�I  jL2  �r�I  h h(h
c__builtin__
__main__
hNN}r�I  Ntr�I  Rr�I  �r�I  Rr�I  X   NNr�I  G?�      sX   RBSr�I  jb  �r�I  h h(h
c__builtin__
__main__
hNN}r�I  Ntr�I  Rr�I  �r�I  Rr�I  X   JJr�I  G?�      sX   JJSr�I  j  �r�I  h h(h
c__builtin__
__main__
hNN}r�I  Ntr�I  Rr�I  �r�I  Rr�I  X   NNr�I  G?�      sX   ``r�I  j�<  �r�I  h h(h
c__builtin__
__main__
hNN}r�I  Ntr�I  Rr�I  �r�I  Rr�I  X   VBZr�I  G?�      su.