�cdill._dill
_load_type
q X   setq�qRq]q(X   JJqX   VBZqX   VBPqX   DTqX   JJRq	X   VBq
X   WDTqX   ``qX   VBGqX   NNSqX   RBSqX   CCqX   RBqX   CDqX   NNPSqX   MDqX   PRPqX   .qX   ,qX   WPqX   VBNqX   RPqX   POSqX   oovqX   NNqX   JJSqX   VBDqX   TOq X   INq!X   NNPq"X   ''q#X   WRBq$X   PRP$q%e�q&Rq'.